library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity img_rom is
   port(
      clock         : in std_logic;

      line_data     : in std_logic_vector(10 downto 0);
      column_data   : in std_logic_vector(10 downto 0);

      frst_pixel_h  : in std_logic_vector(10 downto 0);
      frst_pixel_v  : in std_logic_vector(10 downto 0);

      data          : out std_logic_vector(23 downto 0)
		);
end img_rom;

architecture Behavioral of img_rom is
   signal tx: std_logic_vector(23 downto 0);
   type rom_type is array(0 to 159, 0 to 329) of std_logic_vector(23 downto 0);
   
   -- ROM definition
constant ROM: rom_type :=(
(X"FEFFFF",X"D7D6D2",X"FFC1AD",X"FFACBF",X"FFA2B0",X"FFABAE",X"FFACAF",X"FF9EAE",X"FFA2B2",X"FFAEB4",X"FFAAB8",X"FFAABA",X"FFB2C4",X"E7CFCF",X"D8D6D7",X"BCD9D4",X"7AFFE2",X"8EFFF8",X"8AFFF7",X"7CFFF6",X"82FFF6",X"7BFFF3",X"76FFF4",X"99F6EE",X"CFD9D1",X"E2C8D1",X"FFC4E9",X"FF9CDE",X"FF9FEC",X"FFA7F3",X"FF97E8",X"FF9BE3",X"FF9BE5",X"FFA5F3",X"FFBBD8",X"E2D0CE",X"C8D2F6",X"ADE1FF",X"9DF2FF",X"99E2FF",X"A8E5FF",X"BFD2F3",X"D0CFD5",X"ECD1E2",X"FFB1EE",X"FF9AEB",X"FFA4F1",X"FF9EE8",X"FF9CF4",X"FF91EF",X"FFA4F6",X"FFBDE9",X"E3CACE",X"D3D5D2",X"B8DCEA",X"A4EEFF",X"96E8FF",X"93E9FF",X"9AEEFF",X"9DE4FF",X"ABE7FF",X"A3DEFF",X"9FE4FF",X"99E7FF",X"91E8FF",X"93E8FF",X"95E6FF",X"9CEAFF",X"9BE7FF",X"98E2FF",X"9DE7FF",X"97E3FF",X"9DE9FF",X"9AE6FF",X"98E7FF",X"98E7FF",X"99E4FF",X"9FE6FF",X"A3E4FF",X"9FDFFF",X"A4E3FF",X"99EBFF",X"99ECFF",X"A1E1FF",X"A2E5FF",X"9AE9FF",X"A4E2FF",X"CBE3FF",X"CFD8D7",X"CED1DA",X"DFD6EB",X"D7D1DD",X"DCCFBF",X"FFC6A6",X"FFCE84",X"FFD178",X"FFCA72",X"FFCF68",X"FFCE70",X"FFC891",X"FFCEAE",X"D5D0D4",X"E1D5E3",X"C2E0BC",X"CFFEC7",X"CAEEC0",X"D8EBCB",X"ECF0DF",X"FFFEFA",X"FDF7F9",X"F9F6FD",X"FEFEFF",X"FFFFF8",X"FDF2FF",X"FFFDFF",X"F9FFF6",X"FDFCF7",X"F6E3DC",X"DCD2C8",X"CBD6DA",X"C8D4FF",X"A6DEFF",X"A0EAFF",X"9EE0FF",X"96E4FF",X"98E1FF",X"A5E6FF",X"9DE1FF",X"A0E5FF",X"E0F7FF",X"FFF8F7",X"FFFBFF",X"F3FEFF",X"F6FBFE",X"FFFEFF",X"FCF5FD",X"C2DDF2",X"CAC9FF",X"AAE4FF",X"99EEFF",X"95DDFF",X"9CEAFF",X"A5EBFF",X"8AE4FF",X"ABE7FF",X"B8D8FF",X"D2D9E3",X"F5F6EE",X"F5FAFE",X"FAF6ED",X"FFD5BA",X"FFC668",X"FFC871",X"FFD46F",X"FFCC7E",X"FFCB89",X"FFC599",X"CDCED0",X"D7DCF0",X"D0E8C6",X"D0F5B0",X"E0FDC5",X"F0FFED",X"F9FEFF",X"FFFCFF",X"F8F8F6",X"F8FCFB",X"FFFBFF",X"FDFDFF",X"FEFEFF",X"FFFFFF",X"FFFFFD",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FDFEFF",X"FFFAF8",X"F6FDF5",X"FAFFFA",X"FFFBFF",X"FFFDFF",X"F2F7FD",X"D5FFFF",X"90FFE8",X"8DFFEF",X"96FAF0",X"B7F0E9",X"CED9D1",X"DAD0E8",X"BCCFFF",X"A6E2FF",X"9FE7FF",X"8FE9FF",X"A0E5FF",X"AFD7FF",X"CCDAF7",X"FFF9FF",X"FFF9FD",X"FFFFFB",X"F6FFF8",X"DAD5D2",X"F0F275",X"FFFF6A",X"FFF66C",X"FFF36C",X"FFF9AA",X"E3E1CA",X"CDD0D5",X"D7CCDA",X"F2C4CF",X"FFB4E2",X"FCF1ED",X"F8FFFF",X"F8FEFA",X"FFFEFF",X"FFFFFB",X"FDFFFE",X"FFF7FA",X"FFFFFF",X"FAFBFF",X"F9F9FF",X"C9E9E8",X"C2EAE9",X"D8D7E5",X"D5D0D7",X"F0C3E0",X"FFB1EA",X"FF9FE8",X"FFA9ED",X"FFB4E2",X"ECCBE0",X"D7D2D6",X"C4DDFF",X"A5DBFF",X"A2E0FF",X"ACDDFF",X"A8DBFF",X"AAE8FF",X"B3D4FF",X"E2D2DC",X"DACBD2",X"FFB2EC",X"FFA2EE",X"FFA8E1",X"FFA8E1",X"FFA0EF",X"FFA2F4",X"FFA2EC",X"FFA5E9",X"FFA9EC",X"FFA4E9",X"FFA0ED",X"FFA1EF",X"FFACF2",X"FFA9EC",X"FFA9ED",X"E5CEE8",X"E6D1E4",X"D5C8D1",X"D8DDD7",X"C2D9C7",X"B8DAC1",X"C5E3C9",X"C2DAC2",X"DAD3DA",X"BEE0D0",X"D9D7C8",X"FFCFB4",X"FFC380",X"FFD56B",X"FFD77F",X"FFCE98",X"D6D5C3",X"D1D2CD",X"E0E6A8",X"F5F281",X"F9E07C",X"FFE97B",X"FFEB65",X"FFEE7B",X"FFE96A",X"FBEB72",X"FFEC76",X"FFE97A",X"F4DC92",X"D1D5C6",X"EAD7F7",X"FFBDF3",X"FFA5EE",X"FFA4ED",X"FFC2EF",X"DECCCC",X"CED1C8",X"DBDAE2",X"C1DFE7",X"A4FAED",X"80FDF7",X"8FFFFF",X"8BFFF0",X"95FEED",X"95FAE8",X"97FFF0",X"95FFF5",X"8BFFF2",X"B3E0DD",X"C2E2E1",X"CBD9DC",X"DBCFDB",X"F2C7E3",X"FFBCEC",X"FFA2E8",X"FFA2F6",X"FFABEF",X"FFA3F1",X"FFA3F6",X"FFA8F5",X"FFB4F2",X"FFACE3",X"FFA5E3",X"FFB1F8",X"D6D1E5",X"D5CBD4",X"D6D6D8",X"C5E2EA",X"ABE2FF",X"9EE1FF",X"9FE5FF",X"9EEAFF",X"AEDCFF",X"F1EFFF"),
(X"FEFFFF",X"858480",X"4D0000",X"7D081B",X"8C000C",X"841114",X"7A0D10",X"940B1B",X"8F0111",X"780D13",X"850816",X"780818",X"5E000D",X"180000",X"010000",X"001712",X"199E81",X"209F8A",X"239D90",X"17A491",X"139E87",X"12A78A",X"13B091",X"126F67",X"000400",X"150004",X"48001D",X"940F51",X"8D0D5A",X"86105C",X"9D0B5C",X"9F175F",X"91115B",X"8F1260",X"450019",X"0F0000",X"00092D",X"114581",X"055A91",X"1760A4",X"0A4786",X"000526",X"05040A",X"110007",X"61013E",X"951061",X"8A0B58",X"90125C",X"9B0C64",X"A10C6A",X"8E1062",X"4D0632",X"130000",X"000100",X"001B29",X"095370",X"14669E",X"0E6493",X"085C8B",X"0B5290",X"14508F",X"1E5991",X"185D98",X"0B59A1",X"075EA1",X"1267A7",X"1566A5",X"12609E",X"0E5A98",X"135D9C",X"17619E",X"09558F",X"07538F",X"05518B",X"0B5A92",X"12619A",X"105B9C",X"0D5496",X"105193",X"11518F",X"165598",X"0A5C8C",X"156894",X"185895",X"0A4D94",X"025193",X"135180",X"000327",X"000302",X"00030C",X"040010",X"08020E",X"0C0000",X"8D3A1A",X"C38339",X"BE741B",X"CC7820",X"C57C15",X"C07E20",X"D0753E",X"744323",X"030002",X"070009",X"375531",X"77A66F",X"94B88A",X"8B9E7E",X"E5E9D8",X"FFFAF6",X"FEF8FA",X"FFFDFF",X"FEFEFF",X"FAFAF2",X"FFF8FF",X"FCF7FD",X"FBFFF8",X"FBFAF5",X"A18E87",X"0D0300",X"000408",X"000B53",X"0A4295",X"004778",X"1D5F8F",X"115F90",X"054E9B",X"1B5C9C",X"094D96",X"135881",X"C3DAEA",X"FFFCFB",X"FAF5F9",X"F3FEFF",X"F9FEFF",X"FFFDFE",X"F3ECF4",X"001126",X"03023E",X"0A4483",X"065B91",X"0A528C",X"0C5A9A",X"084E93",X"0B659A",X"235F91",X"000536",X"00010B",X"ECEDE5",X"FBFFFF",X"FEFAF1",X"D3A186",X"C46B0D",X"CD6D16",X"AE7A15",X"B96C1E",X"C97836",X"6C2C00",X"020305",X"000013",X"6E8664",X"7EA35E",X"84A169",X"D3E6D0",X"FBFFFF",X"FEF9FF",X"FEFEFC",X"FCFFFF",X"FFFDFF",X"FDFDFF",X"FEFEFF",X"FFFFFF",X"FFFFFD",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FDFEFF",X"FFF2F0",X"FBFFFA",X"F7FEF7",X"FFF5F9",X"FEFCFF",X"FAFFFF",X"C9FCF5",X"198E71",X"19987B",X"35998F",X"0B443D",X"000400",X"040012",X"000C4E",X"134F95",X"0D5587",X"0B6599",X"02478C",X"00215E",X"98A6C3",X"FFFAFF",X"FFF6FA",X"FFFFFB",X"EAF4EC",X"140F0C",X"BCBE41",X"DFD540",X"E2CB41",X"E6D24B",X"C0B566",X"040200",X"04070C",X"07000A",X"2C0009",X"69103E",X"E7DCD8",X"F8FFFF",X"FAFFFC",X"FCFAFF",X"FFFFFB",X"FEFFFF",X"FFF6F9",X"FBFBFD",X"FEFFFF",X"FBFBFF",X"739392",X"012928",X"00000C",X"030005",X"390C29",X"63013A",X"8D0F58",X"840F53",X"520533",X"17000B",X"030002",X"051E60",X"104684",X"094782",X"18498C",X"003081",X"0F4D98",X"001845",X"0A0004",X"14050C",X"66013B",X"890652",X"7F124B",X"84114A",X"880958",X"80095B",X"830B55",X"860F53",X"7C0F52",X"811257",X"90105D",X"870A58",X"751056",X"670649",X"6F0448",X"0E0011",X"0D000B",X"0B0007",X"000200",X"001100",X"12341B",X"5A785E",X"5C745C",X"040004",X"000E00",X"0D0B00",X"AF6F54",X"E18A47",X"BF8016",X"BB7B23",X"9B5E28",X"0A0900",X"000100",X"42480A",X"A9A635",X"B9A03C",X"B49022",X"C4A21C",X"C6A532",X"B8991A",X"B1A128",X"B29923",X"C69E2F",X"826A20",X"000300",X"2F1C3C",X"6B255B",X"860A53",X"8D135C",X"540532",X"150303",X"010400",X"010008",X"001B23",X"277D70",X"08857F",X"179389",X"168B7B",X"0F7867",X"1F8472",X"299482",X"0E7E6E",X"188C7F",X"13403D",X"000C0B",X"000407",X"080008",X"280019",X"590B3B",X"810F55",X"860052",X"8B1458",X"850856",X"8D0C5F",X"7D0350",X"952967",X"7B184F",X"7A1654",X"6C054C",X"010010",X"0D030C",X"000002",X"000810",X"245B7A",X"105387",X"00427D",X"0D598D",X"001450",X"CECCF4"),
(X"FFF0FB",X"BE828E",X"900000",X"D43150",X"D61B36",X"D21A32",X"CA122E",X"D21535",X"D31C38",X"D21B39",X"DF153D",X"C12645",X"6C242F",X"261C1B",X"021010",X"377568",X"1FC7A3",X"1CC5A4",X"1DC1A8",X"14C7A9",X"17C2A2",X"16BF9E",X"24CDAC",X"1C867C",X"10060F",X"191C23",X"7C1A4D",X"E92D8C",X"EC1187",X"ED0C8C",X"D7168B",X"DE178B",X"CF1B7E",X"9C306E",X"3A1830",X"000E33",X"215CAC",X"2387DC",X"0D7BD2",X"1272EA",X"1D7DEB",X"2A60C4",X"002556",X"102422",X"4F212B",X"AB3572",X"DE2791",X"FB0B88",X"F1147B",X"EC1A85",X"DE1D88",X"C71A76",X"9C1758",X"520732",X"200C2F",X"29375A",X"4578BA",X"3A7CC8",X"267EE0",X"1E8DFF",X"0C8BFC",X"0A8CEA",X"067FDC",X"0C78E4",X"117FF2",X"0F7EEA",X"0D7DDF",X"1381E2",X"107EE0",X"117CE4",X"1D88F2",X"208BF5",X"147CEB",X"1379E5",X"187AE5",X"1B7BE9",X"1675E9",X"1472EE",X"1776F6",X"187AF9",X"1C8AFD",X"0B74E9",X"137DEA",X"1D80DD",X"377FC9",X"406496",X"24344E",X"03111C",X"000600",X"080300",X"2D2226",X"1E1B24",X"1C1000",X"C6693D",X"EB8A29",X"F98410",X"FF7C1F",X"FD7E0D",X"F37E15",X"FD823C",X"9A572C",X"130900",X"130907",X"748F58",X"85AE72",X"89A87C",X"BACAB0",X"FAFBF6",X"FFFCFF",X"FFFAFF",X"FCFAFD",X"FDFFFC",X"FFFDFA",X"F7FDFB",X"F6FFFF",X"FFF0E0",X"FFD39A",X"C46D38",X"5C1A0E",X"1D040A",X"2C2C46",X"3F78AF",X"1B81E6",X"0E74D6",X"2076E7",X"1B7FE1",X"1480E2",X"076EB3",X"88B5D2",X"F7FFFF",X"FFFAFA",X"F9F3F5",X"FCFFFF",X"F7F9F6",X"F9F9F7",X"F0F5FB",X"4079C0",X"2C61CB",X"247FF2",X"1284E7",X"117FE1",X"1B81F0",X"1574E0",X"1F83D9",X"3F6E9A",X"243455",X"070000",X"E7D9CE",X"FFFFFF",X"F5F6F1",X"FFE9DB",X"C18A4A",X"F77227",X"FA7B12",X"FF7A1A",X"F1763A",X"82412D",X"1A1617",X"0F1E0B",X"6F9D55",X"86B871",X"88B270",X"9FBB93",X"ECF7EF",X"FBF9FE",X"FFFFFD",X"F0F2ED",X"FCFCFE",X"FDFCFF",X"FEFEFF",X"FFFFFF",X"FFFFFD",X"FFFFFD",X"FFFFFF",X"FEFFFF",X"FDFEFF",X"F5FFFF",X"F5F8FD",X"FFFCFF",X"FAFFFE",X"FEF8FC",X"E4FFFF",X"79DAC7",X"09AF8B",X"29AC9A",X"449C90",X"202F34",X"0F0D22",X"0C3B69",X"246EC7",X"1E69DC",X"1270E1",X"1C6FE9",X"2A69CA",X"577AB4",X"DFECFC",X"FFFFF8",X"FFFAFA",X"FFFEFD",X"EAECD7",X"91883D",X"E0E121",X"E3D804",X"F1D51C",X"E9D542",X"696827",X"000400",X"292E32",X"441120",X"AC2462",X"BB006A",X"FFD1F3",X"FEFFFF",X"FFFFF1",X"FFF9FF",X"F6FFFF",X"FFF9FF",X"FFFDFB",X"FCFFFB",X"F5FFFF",X"E5F6F0",X"536A58",X"000300",X"3E1F25",X"4A0035",X"99276D",X"DE3E98",X"D71B7C",X"CA2076",X"901F55",X"3F1628",X"111811",X"134286",X"2977DB",X"1979EA",X"156DD1",X"1569C9",X"3184E2",X"26589D",X"121737",X"2F1A2D",X"8F1D62",X"CA1F85",X"CE1A7E",X"D61679",X"DB187E",X"D91C83",X"E41F89",X"CD0F71",X"D11979",X"CD2079",X"BF2875",X"9A2D66",X"7D3D5F",X"5C3748",X"3B1B26",X"152115",X"283B28",X"355138",X"547C59",X"6B986F",X"77A87B",X"84B888",X"84B888",X"4E5840",X"231316",X"0E0004",X"A05D4C",X"F49658",X"F97F2C",X"DD7B22",X"FB8B43",X"743514",X"290914",X"3A3434",X"9D9445",X"E3C23D",X"CDA61B",X"C2AC18",X"BFBC0F",X"D8B71C",X"B49F06",X"C9B018",X"CDAA1C",X"CCB545",X"65622B",X"13000B",X"6C356F",X"AF3D92",X"CE2693",X"D9228E",X"9F1D63",X"500E34",X"2D0C2B",X"050414",X"41625B",X"50968B",X"1E9881",X"009F81",X"21BDA7",X"21B4A4",X"0EA997",X"0FAE9A",X"0FA896",X"31A495",X"228378",X"003431",X"35535D",X"3E344D",X"713B6C",X"973A80",X"9F2A7B",X"AB095C",X"C4247E",X"BA1679",X"D3298C",X"BB0C6B",X"CC1774",X"D01B7A",X"E83296",X"A81D6E",X"6D194D",X"2F0D2E",X"22173F",X"414A8B",X"3664BA",X"1A64C7",X"2879E4",X"0051A1",X"BEE4FF"),
(X"FFF2FD",X"CA8E9A",X"9C0806",X"C52241",X"C50A25",X"C00820",X"C8102C",X"C70A2A",X"C00925",X"BF0826",X"CC022A",X"AD1231",X"4E0611",X"0A0000",X"061414",X"559386",X"1BC39F",X"1BC4A3",X"12B69D",X"08BB9D",X"18C3A3",X"07B08F",X"1BC4A3",X"309A90",X"080007",X"000007",X"741245",X"CE1271",X"DC0177",X"E50484",X"CD0C81",X"D40D81",X"D52184",X"7D114F",X"1D0013",X"010F34",X"2F6ABA",X"177BD0",X"0D7BD2",X"0B6BE3",X"0E6EDC",X"3268CC",X"295182",X"051917",X"240000",X"800A47",X"C60F79",X"F0007D",X"E3066D",X"D90772",X"CB0A75",X"C61975",X"AF2A6B",X"6A1F4A",X"180427",X"000023",X"001355",X"1E60AC",X"277FE1",X"0D7CF2",X"0483F4",X"0A8CEA",X"0780DD",X"1581ED",X"117FF2",X"0675E1",X"0070D2",X"0A78D9",X"0775D7",X"016CD4",X"0C77E1",X"147FE9",X"0B73E2",X"0C72DE",X"0F71DC",X"0E6EDC",X"0C6BDF",X"1270EC",X"1675F5",X"1173F2",X"0573E6",X"1D86FB",X"0A74E1",X"187BD8",X"1860AA",X"05295B",X"00021C",X"14222D",X"717755",X"625D4A",X"070000",X"09060F",X"1A0E00",X"D27549",X"E68524",X"ED7804",X"FF7417",X"FD7E0D",X"F37E15",X"F27731",X"844116",X"080000",X"090000",X"76915A",X"87B074",X"77966A",X"E9F9DF",X"F7F8F3",X"FDF6FD",X"FEF7FF",X"FBF9FC",X"FEFFFD",X"FFFBF8",X"F3F9F7",X"F7FFFF",X"FFF2E2",X"F0B37A",X"CC7540",X"A46256",X"130000",X"090923",X"1A538A",X"076DD2",X"0C72D4",X"1066D7",X"1377D9",X"107CDE",X"0970B5",X"BBE8FF",X"F7FFFF",X"FFF3F3",X"FCF6F8",X"FCFFFF",X"FDFFFC",X"FFFFFD",X"E8EDF3",X"427BC2",X"285DC7",X"0A65D8",X"0577DA",X"0775D7",X"0A70DF",X"1E7DE9",X"1377CD",X"174672",X"000122",X"0C0300",X"F4E6DB",X"FCFCFE",X"FAFBF6",X"FFF1E3",X"FDC686",X"E96419",X"F2730A",X"FF6B0B",X"EF7438",X"7B3A26",X"1D191A",X"172613",X"719F57",X"7BAD66",X"85AF6D",X"84A078",X"B4BFB7",X"FFFEFF",X"F7F6F4",X"FEFFFB",X"FEFEFF",X"FDFCFF",X"FEFEFF",X"FFFFFF",X"FFFFFD",X"FFFFFD",X"FFFFFF",X"FEFFFF",X"FDFEFF",X"F4FFFF",X"FCFFFF",X"FFFAFF",X"F7FDFB",X"FFFDFF",X"D7FAF6",X"4BAC99",X"17BD99",X"2DB09E",X"004B3F",X"000409",X"010014",X"31608E",X"2973CC",X"1863D6",X"116FE0",X"176AE4",X"1554B5",X"A6C9FF",X"F4FFFF",X"F8F8F0",X"FAF4F4",X"FAF6F5",X"F8FAE5",X"C9C075",X"E3E424",X"EFE410",X"FBDF26",X"E5D13E",X"474605",X"020A00",X"12171B",X"410E1D",X"B62E6C",X"C0006F",X"FFCDEF",X"FEFFFF",X"F5F6E6",X"FFF9FF",X"F7FFFF",X"FFFCFF",X"FFF9F7",X"F5FAF4",X"F3FFFF",X"F3FFFE",X"5C7361",X"000200",X"47282E",X"6F225A",X"98266C",X"E4449E",X"CD1172",X"C51B71",X"8D1C52",X"2F0618",X"020902",X"09387C",X"1A68CC",X"0C6CDD",X"035BBF",X"166ACA",X"1E71CF",X"23559A",X"0B1030",X"130011",X"760449",X"BA0F75",X"C10D71",X"C8086B",X"CB086E",X"C1046B",X"C7026C",X"D11375",X"BB0363",X"BC0F68",X"A10A57",X"680034",X"360018",X"180004",X"180003",X"414D41",X"708370",X"7D9980",X"87AF8C",X"74A178",X"5E8F62",X"598D5D",X"76AA7A",X"727C64",X"0B0000",X"0F0005",X"8A4736",X"DD7F41",X"F47A27",X"E17F26",X"F08038",X"B87958",X"1C0007",X"040000",X"605708",X"CFAE29",X"CEA71C",X"C1AB17",X"C5C215",X"CCAB10",X"B9A40B",X"CCB31B",X"D6B325",X"C8B141",X"8A8750",X"0D0005",X"69326C",X"9A287D",X"B60E7B",X"C30C78",X"AB296F",X"5E1C42",X"2E0D2C",X"00000F",X"000C05",X"1C6257",X"26A089",X"07A688",X"12AE98",X"16A999",X"0EA997",X"18B7A3",X"10A997",X"39AC9D",X"49AA9F",X"3C817E",X"2F4D57",X"060015",X"34002F",X"7D2066",X"931E6F",X"D53386",X"B81872",X"AF0B6E",X"B80E71",X"E03190",X"C81370",X"D01B7A",X"BA0468",X"A4196A",X"B15D91",X"6E4C6D",X"0B0028",X"000243",X"305EB4",X"2973D6",X"1465D0",X"0053A3",X"AED4FF"),
(X"FFFDFD",X"D87B8D",X"BD0000",X"CE1736",X"D10A27",X"DB0024",X"E10027",X"D40026",X"CF0326",X"DD002A",X"E90030",X"B51032",X"270E0A",X"000400",X"0C3B35",X"36B799",X"0DCAA2",X"07CEA7",X"02C1A2",X"00C3A1",X"0ACEAA",X"00BB95",X"14CEA9",X"2CB1A0",X"18272A",X"06050D",X"661840",X"CC1A70",X"DD0B79",X"D40780",X"D90283",X"DF0A8A",X"A61A71",X"2E042A",X"000607",X"295272",X"2876DB",X"056AF6",X"0F71F6",X"0569E1",X"056CEC",X"1875F6",X"1F71DF",X"07387D",X"010017",X"33010D",X"7F224E",X"BB2C86",X"C50D7D",X"E90985",X"F30581",X"DB0778",X"CF0F76",X"CC1476",X"9C0E62",X"570040",X"190007",X"0A0313",X"2D4F74",X"3F82C9",X"237AD7",X"1C7DDB",X"288CEC",X"0C71D9",X"137CEF",X"1180EC",X"0A7DEA",X"077CF0",X"0176F7",X"0477F8",X"0B7EF3",X"0378E1",X"0473E9",X"0273E9",X"087AEC",X"097DEC",X"037AE2",X"0077D8",X"0078D3",X"0078CE",X"1772CF",X"307ED1",X"5483C9",X"303869",X"040015",X"160C15",X"080004",X"4D3C46",X"D9D4B6",X"C2B299",X"070000",X"15161B",X"120600",X"DC7942",X"F77F0F",X"FF7E00",X"F47504",X"F57B00",X"FA8406",X"F7862A",X"7C460A",X"010200",X"080E02",X"879F63",X"91AF79",X"AEC49E",X"F7FFF2",X"FFFDFF",X"FBF2FF",X"FFFBFF",X"FEFEFE",X"F7FAF1",X"FCF7FE",X"F7FFFF",X"F6F3EE",X"FFDBB4",X"F67E1D",X"FB780C",X"DE7B37",X"602500",X"020403",X"05000D",X"375392",X"2378B9",X"0C6DD4",X"1276F0",X"055CC6",X"76B0C8",X"EEFCFF",X"FFFEFF",X"FFFBFB",X"FFFBFC",X"F6F2EF",X"FEFEF6",X"FBFFFD",X"E4F5FC",X"3983D8",X"046CDF",X"0777F7",X"118AF3",X"067FDC",X"0A6BD6",X"2B7CD8",X"2369A5",X"041028",X"110101",X"381300",X"FBDCCA",X"FFFDFF",X"F9FFFF",X"FCF8F5",X"FFEED8",X"E09159",X"EC720D",X"FF7600",X"E06B28",X"4E2C2A",X"070105",X"1B3005",X"7EB365",X"71AF64",X"7CB566",X"7CA364",X"3C4E34",X"E9EAEC",X"FAF4F4",X"FFFCF7",X"FBFFFF",X"FEFCFF",X"FFFDFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FDFEFF",X"FFFBFA",X"FFFAFD",X"F7FFFF",X"F5F6FB",X"E4FFFF",X"8CE9DE",X"02A68B",X"1FB09F",X"2B7F6F",X"000A18",X"00022C",X"034083",X"2276D6",X"0064D3",X"0069E1",X"1268EF",X"175FE5",X"366BB9",X"D4ECFF",X"F7FFFF",X"FCFFF1",X"FEFFFF",X"FCF6F6",X"FFFDCB",X"F4E25C",X"E2D400",X"EADA0B",X"E1D146",X"AFA756",X"0D0000",X"180A0A",X"211215",X"1B0709",X"861D56",X"B20E6D",X"FFD2EF",X"F8FBFF",X"FFFCFB",X"FFFAFF",X"EDF9EF",X"FDFDFF",X"FAFDF2",X"FFFFFA",X"FCFAFF",X"FBEDFF",X"995A77",X"6A0025",X"B31C6B",X"C3127C",X"C20271",X"D40075",X"D5006D",X"CF046F",X"B62777",X"4D0B39",X"040012",X"19294B",X"295EBC",X"1065E4",X"0B67D4",X"116ECD",X"136ED7",X"165BBA",X"0A3071",X"00050F",X"490735",X"A51368",X"CB0B7C",X"D70075",X"D7066E",X"CD026E",X"DA007B",X"BB0063",X"C11A76",X"710042",X"2A001B",X"010302",X"001500",X"4F7D4E",X"609A5F",X"6EA56B",X"6DAB6C",X"6CAF6C",X"5D9B58",X"629958",X"649254",X"709E60",X"649456",X"70A169",X"404C36",X"0D0000",X"363022",X"CB7954",X"ED7E2F",X"FF801E",X"F47D15",X"F2863D",X"9B512C",X"170000",X"0F0500",X"8A7A25",X"D5B52C",X"C2A605",X"BDB009",X"CCA605",X"DEBD16",X"C1A000",X"C5A502",X"D9C028",X"B7A539",X"180200",X"735587",X"A54585",X"A0086D",X"C6047E",X"C20470",X"B30A65",X"A71566",X"56002D",X"1B0004",X"0D0000",X"214E47",X"2F978C",X"28AAA0",X"0EAB9A",X"06BD9F",X"07B194",X"23A895",X"05A38C",X"1AA892",X"31A290",X"4A9C8E",X"053831",X"00080B",X"3E3645",X"1C0319",X"7B4263",X"8A2865",X"AC1677",X"BE077D",X"D2158D",X"B10066",X"D11880",X"D7187F",X"BD007B",X"C81D8D",X"AD3889",X"3D083E",X"0B002A",X"1D1F5A",X"305198",X"2C70BB",X"074AB2",X"BFDFFF"),
(X"FFFAFA",X"DF8294",X"CB060D",X"D92241",X"CB0421",X"DE0027",X"DF0025",X"DF0831",X"CE0225",X"DD002A",X"E90030",X"B00B2D",X"1C0300",X"000400",X"1B4A44",X"36B799",X"0CC9A1",X"00C69F",X"05C4A5",X"00C7A5",X"04C8A4",X"07C49E",X"16D0AB",X"21A695",X"000A0D",X"000007",X"52042C",X"CC1A70",X"DB0977",X"D0037C",X"E0098A",X"DF0A8A",X"8C0057",X"280024",X"000607",X"285171",X"3381E6",X"066BF7",X"0B6DF2",X"1175ED",X"0A71F1",X"0A67E8",X"2577E5",X"2F60A5",X"0F0925",X"220000",X"470016",X"A71872",X"CA1282",X"E40480",X"EB0079",X"DA0677",X"CC0C73",X"CF1779",X"B6287C",X"82296B",X"240212",X"03000C",X"001237",X"00357C",X"0F66C3",X"1E7FDD",X"2589E9",X"167BE3",X"137CEF",X"0E7DE9",X"077AE7",X"077CF0",X"0277F8",X"0477F8",X"0C7FF4",X"087DE6",X"0978EE",X"0070E6",X"0375E7",X"0A7EED",X"047BE3",X"0076D7",X"057ED9",X"108AE0",X"1F7AD7",X"0E5CAF",X"103F85",X"000233",X"040015",X"130912",X"0D0409",X"100009",X"8E896B",X"8C7C63",X"070000",X"0F1015",X"100400",X"C15E27",X"FF8E1E",X"FC7100",X"FF800F",X"F97F00",X"FA8406",X"F68529",X"804A0E",X"050600",X"181E12",X"88A064",X"83A16B",X"D2E8C2",X"F6FEF1",X"FFFDFF",X"FFF9FF",X"FFFCFF",X"FCFCFC",X"FEFFF8",X"FBF6FD",X"F6FFFF",X"FFFEF9",X"F6B891",X"E46C0B",X"FE7B0F",X"E6833F",X"965B2F",X"000100",X"0E0516",X"001554",X"1166A7",X"0E6FD6",X"0D71EB",X"085FC9",X"B9F3FF",X"F4FFFF",X"F5F3F8",X"FFF4F4",X"FFFCFD",X"FFFEFB",X"FFFFF8",X"F2F8F4",X"E7F8FF",X"3A84D9",X"0066D9",X"0A7AFA",X"037CE5",X"057EDB",X"1D7EE9",X"1F70CC",X"004480",X"00051D",X"0F0000",X"957046",X"FFEAD8",X"FFF9FB",X"F3FCF9",X"FFFDFA",X"FFFCE6",X"FFC78F",X"DD6300",X"FF7E04",X"D25D1A",X"2F0D0B",X"080206",X"465B30",X"7EB365",X"76B469",X"659E4F",X"9AC182",X"0B1D03",X"A1A2A4",X"FFFDFD",X"FFFEF9",X"F6FBFF",X"FEFCFF",X"FFFDFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FDFEFF",X"FFFEFD",X"FAEBEE",X"F7FFFF",X"FDFEFF",X"D6FDFC",X"57B4A9",X"06AA8F",X"1DAE9D",X"004131",X"000513",X"11244E",X"2D6AAD",X"0A5EBE",X"066CDB",X"0068E0",X"1C72F9",X"0044CA",X"8BC0FF",X"EAFFFF",X"F5FDFF",X"F7FEEC",X"FBFCFE",X"FFFDFD",X"FCF6C4",X"E3D14B",X"EADC00",X"F0E011",X"CDBD32",X"2E2600",X"110400",X"0A0000",X"0A0000",X"281416",X"700740",X"9E0059",X"FFDEFB",X"FBFEFF",X"FDF9F8",X"FFF7FF",X"F8FFFA",X"FFFFFF",X"F9FCF1",X"FDFCF7",X"FBF9FF",X"FAECFF",X"AC6D8A",X"8A0F45",X"BE2776",X"BC0B75",X"CE0E7D",X"D20073",X"DE0076",X"D30873",X"B62777",X"712F5D",X"0E041C",X"000628",X"1247A5",X"0F64E3",X"0662CF",X"106DCC",X"0A65CE",X"2065C4",X"264C8D",X"000913",X"380024",X"960459",X"C70778",X"D20070",X"D20169",X"D00571",X"E30984",X"CC0B74",X"B8116D",X"841355",X"1D000E",X"454746",X"90AD91",X"8FBD8E",X"6EA86D",X"5E955B",X"5F9D5E",X"5C9F5C",X"5C9A57",X"689F5E",X"6F9D5F",X"6F9D5F",X"6C9C5E",X"6D9E66",X"636F59",X"0E0001",X"120C00",X"984621",X"F08132",X"FF8826",X"EB740C",X"FC9047",X"C97F5A",X"2B0C07",X"0A0000",X"4F3F00",X"C4A41B",X"D1B514",X"B9AC05",X"D4AE0D",X"D0AF08",X"DDBC15",X"C9A906",X"C4AB13",X"B8A63A",X"250F00",X"47295B",X"AF4F8F",X"B0187D",X"BC0074",X"C70975",X"B80F6A",X"A61465",X"812358",X"2A0113",X"0E0000",X"00110A",X"00655A",X"37B9AF",X"22BFAE",X"00B294",X"00A386",X"1BA08D",X"0EAC95",X"27B59F",X"219280",X"429486",X"5B8E87",X"384D50",X"06000D",X"0F000C",X"2C0014",X"72104D",X"AA1475",X"EB34AA",X"CB0E86",X"CC1281",X"CC137B",X"E2238A",X"C20180",X"B30878",X"9F2A7B",X"541F55",X"0E002D",X"050742",X"0E2F76",X"2468B3",X"0144AC",X"B4D4FF"),
(X"F0FDF4",X"E38691",X"CF0001",X"D81B37",X"C2021B",X"DF042A",X"DF0027",X"D5032A",X"D60429",X"D80027",X"D8002A",X"AA0527",X"0A0000",X"000202",X"044038",X"13B993",X"13C8A5",X"00C7A3",X"06C3A7",X"01C2A5",X"07C4A4",X"0CC8A5",X"05CCA5",X"13B79E",X"003221",X"000E07",X"27101A",X"902251",X"C21C68",X"D3096C",X"E90A77",X"C0136F",X"3D0014",X"190310",X"02000B",X"121C35",X"356498",X"1D72C5",X"0A71D8",X"0076E4",X"026CE2",X"0076EB",X"007BF6",X"1377F1",X"1F59AD",X"000625",X"090715",X"370E30",X"AA2C7D",X"C31F78",X"D80671",X"EC007E",X"F2008D",X"ED008B",X"EB0687",X"E40B7E",X"972062",X"50082D",X"0E0002",X"010302",X"151712",X"18211E",X"203F53",X"356998",X"277DB6",X"2178C7",X"1B78D8",X"1C80E0",X"137DD1",X"0875C7",X"1179D8",X"1478E8",X"1279D6",X"0B71D3",X"0F71D6",X"1975D8",X"2575CE",X"3173BF",X"396EB0",X"3A67A2",X"1D2645",X"070017",X"180013",X"31001D",X"8C125F",X"A91168",X"5C0029",X"1F000B",X"21000F",X"1F0000",X"1A1712",X"05080D",X"150500",X"C3622F",X"F9821C",X"FF8409",X"F4750A",X"FB7E00",X"FC7E03",X"F07D22",X"864712",X"080000",X"131418",X"828864",X"ABBC9A",X"ECF8E0",X"FEFFF8",X"FBF9FE",X"FFFCFF",X"FCF9FF",X"F5F5F7",X"FBFFFA",X"FCFFFF",X"FAF5F1",X"FFE6BB",X"E97E2C",X"FF710B",X"FF8306",X"EF8C0D",X"C76D0D",X"621300",X"250000",X"0A0A0C",X"000D2A",X"435971",X"1F4284",X"7C9ECC",X"FBFFFF",X"FFFEFD",X"FFFEFF",X"FEF9FD",X"F8F4F5",X"FFF8F5",X"FFFEF8",X"FAFFFF",X"E9FBFF",X"357DCF",X"0071D5",X"1175E7",X"1571C4",X"247EBA",X"3667AA",X"233F67",X"040404",X"240000",X"8F4C21",X"C27F30",X"FFE1CC",X"FEF8F8",X"F3FFFF",X"FBFFFF",X"FDFBFC",X"FFF8EB",X"CF9154",X"D47C10",X"D27F3D",X"040000",X"08020E",X"526643",X"8AB482",X"87C876",X"6BAA4F",X"95BE6F",X"546843",X"000104",X"EBDFDF",X"FFFCF6",X"F7FFFF",X"FFFBFF",X"FFFDFF",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FFFFFD",X"FFFFFD",X"FEFEFE",X"FBFCF4",X"FFFCFB",X"FFF1FE",X"E5FFFF",X"9EF1E7",X"06AC88",X"2CA18E",X"173C44",X"000019",X"001046",X"215FB6",X"0D6CD6",X"006CDB",X"0A68D9",X"0D62CD",X"0063C1",X"2D6AA0",X"CBF1FA",X"F0F7FD",X"FFFEFF",X"FCFFF4",X"F2F9FF",X"FFFFFD",X"FFFFBB",X"E5CE42",X"E5D220",X"D8CE5F",X"4C5334",X"070200",X"5B2B27",X"713211",X"945E38",X"070300",X"110708",X"30061A",X"E1E1E3",X"FEFCFF",X"FFFEFF",X"F9F7FF",X"FFFFF2",X"F7FFFF",X"F6FFF3",X"FFFCF7",X"FFF7FF",X"FFE1FF",X"CB5A90",X"BD0259",X"DA1686",X"C70E6C",X"BF176E",X"B31F6D",X"B22A72",X"992360",X"610D3E",X"341330",X"040A18",X"000231",X"0B43A0",X"126CE7",X"0568DD",X"0F74E0",X"0066DB",X"0667DC",X"045AC1",X"00223F",X"050217",X"5F143B",X"B11F70",X"CA0F78",X"CD0A72",X"C80470",X"D10381",X"DE0175",X"BD0567",X"871D5B",X"12000D",X"607564",X"97B089",X"7B9D61",X"5B9145",X"619C4C",X"69A658",X"5A994A",X"5E9E50",X"5C9F52",X"5DA053",X"519548",X"6BAF62",X"5DA565",X"6BA05C",X"27451F",X"000105",X"382A1F",X"DA8243",X"F27B13",X"F38A17",X"E57B0E",X"FA8D3A",X"924B15",X"100200",X"19221F",X"A0974C",X"DAB62A",X"D3A31B",X"C9A10C",X"DFB314",X"D5AD0F",X"CBAA0F",X"D0B00D",X"C7A414",X"553C00",X"04000E",X"5E474F",X"902664",X"C1066F",X"CF016D",X"BB0060",X"C10D71",X"BE1773",X"9D0653",X"2C0013",X"100013",X"00091F",X"275660",X"419B91",X"35B197",X"2DA98F",X"3EA798",X"3F7883",X"386673",X"1D4151",X"001B2E",X"132C42",X"071C37",X"0D2040",X"00082B",X"0C0330",X"1A0435",X"55235E",X"7B1F68",X"AE237C",X"AB0066",X"BE0675",X"B5006D",X"CD006F",X"CD137E",X"B41571",X"981259",X"630134",X"35052B",X"010125",X"364F78",X"144C96",X"B7DCFF"),
(X"F7FFFB",X"E28590",X"CD0000",X"D91C38",X"CA0A23",X"D4001F",X"DF0027",X"D40229",X"D30126",X"D70026",X"D9002B",X"B10C2E",X"0D0000",X"080E0E",X"00372F",X"15BB95",X"12C7A4",X"05CDA9",X"00BDA1",X"00B99C",X"0AC7A7",X"08C4A1",X"00BD96",X"29CDB4",X"3D7C6B",X"000F08",X"160009",X"6E002F",X"CA2470",X"DA1073",X"E50673",X"C11470",X"35000C",X"13000A",X"04020D",X"00031C",X"00194D",X"1C71C4",X"1980E7",X"0076E4",X"0D77ED",X"0077EC",X"007CF7",X"0E72EC",X"3872C6",X"264564",X"00000C",X"1C0015",X"700043",X"B9156E",X"E2107B",X"ED017F",X"F1008C",X"ED008B",X"E90485",X"E2097C",X"9E2769",X"6C2449",X"210C15",X"000201",X"000100",X"000502",X"00091D",X"00204F",X"045A93",X"156CBB",X"1D7ADA",X"1D81E1",X"157FD3",X"1380D2",X"177FDE",X"0C70E0",X"1279D6",X"167CDE",X"197BE0",X"1975D8",X"2373CC",X"2567B3",X"073C7E",X"000A45",X"000928",X"221332",X"3D1538",X"681F54",X"A42A77",X"BD257C",X"8F1E5C",X"4F1E3B",X"421430",X"2F070F",X"090601",X"000005",X"160600",X"D3723F",X"F67F19",X"F47600",X"FB7C11",X"FA7D00",X"F67800",X"FA872C",X"A1622D",X"080000",X"000105",X"656B47",X"D4E5C3",X"F7FFEB",X"F9FCF3",X"FFFEFF",X"FEF8FF",X"FFFCFF",X"FFFFFF",X"F5FAF4",X"F6FAFB",X"FFFBF7",X"F3C89D",X"D66B19",X"FF7C16",X"F97900",X"DF7C00",X"E68C2C",X"C6773C",X"582915",X"000002",X"0B1A37",X"00041C",X"001658",X"C1E3FF",X"FAFEFF",X"FEFAF9",X"FFFCFD",X"FDF8FC",X"FFFEFF",X"FFFDFA",X"FFFBF5",X"FBFFFF",X"DFF1FB",X"357DCF",X"007CE0",X"0C70E2",X"207CCF",X"1E78B4",X"00286B",X"00133B",X"020202",X"532611",X"CA875C",X"BE7B2C",X"FFDAC5",X"FFFDFD",X"F5FFFF",X"F5FBFB",X"FEFCFD",X"FEF6E9",X"FFD295",X"CB7307",X"BB6826",X"040000",X"04000A",X"576B48",X"89B381",X"6BAC5A",X"6DAC51",X"92BB6C",X"617550",X"000306",X"AB9F9F",X"FFFCF6",X"EFF9FF",X"FFFBFF",X"FFFDFF",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FFFFFD",X"FFFFFD",X"FEFEFE",X"FEFFF7",X"FFFBFA",X"FFF5FF",X"DBFDFE",X"79CCC2",X"02A884",X"0C816E",X"001D25",X"00021C",X"25447A",X"2765BC",X"0B6AD4",X"006EDD",X"0361D2",X"1C71DC",X"0062C0",X"72AFE5",X"E0FFFF",X"F8FFFF",X"FEFCFF",X"FBFFF3",X"F7FEFF",X"FFFFFD",X"FEF7B1",X"EDD64A",X"F0DD2B",X"827809",X"050C00",X"130E0B",X"3B0B07",X"C28362",X"C7916B",X"504C29",X"0A0001",X"1B0005",X"E5E5E7",X"FFFEFF",X"FAF9FF",X"FFFDFF",X"FFFFF3",X"F6FFFF",X"F8FFF5",X"FFFAF5",X"FFF7FF",X"FFE2FF",X"C8578D",X"BD0259",X"D71383",X"CF1674",X"BD156C",X"9E0A58",X"8B034B",X"67002E",X"5A0637",X"140010",X"000513",X"0E2352",X"1F57B4",X"035DD8",X"0669DE",X"0061CD",X"066FE4",X"0263D8",X"186ED5",X"0F3C59",X"000012",X"4B0027",X"A21061",X"C20770",X"CA076F",X"C6026E",X"CC007C",X"D6006D",X"C91173",X"821856",X"160011",X"697E6D",X"809972",X"7FA165",X"699F53",X"639E4E",X"5D9A4C",X"65A455",X"5B9B4D",X"5B9E51",X"61A457",X"67AB5E",X"5EA255",X"5FA767",X"6BA05C",X"587650",X"000408",X"0B0000",X"B45C1D",X"F27B13",X"F08714",X"FB9124",X"E87B28",X"D28B55",X"23150A",X"000704",X"6C6318",X"C6A216",X"DDAD25",X"CFA712",X"D7AB0C",X"C59D00",X"DCBB20",X"C9A906",X"CBA818",X"947B38",X"060010",X"19020A",X"9E3472",X"C1066F",X"CD006B",X"C9096E",X"BF0B6F",X"B30C68",X"B01966",X"5F2D46",X"210A24",X"0C172D",X"002C36",X"005A50",X"209C82",X"037F65",X"005D4E",X"002530",X"000E1B",X"000D1D",X"000E21",X"000C22",X"011631",X"031636",X"162447",X"1F1643",X"13002E",X"34023D",X"6E125B",X"A21770",X"B90E74",X"BF0776",X"C00578",X"D40476",X"BE046F",X"CE2F8B",X"BE387F",X"811F52",X"36062C",X"000023",X"0C254E",X"002B75",X"BCE1FF"),
(X"FCFBF7",X"E7838D",X"D50000",X"E51836",X"D00321",X"D70329",X"DC012B",X"DA042A",X"DB0026",X"D00025",X"D60029",X"C70A32",X"310708",X"040000",X"073832",X"2BB79A",X"14CCA6",X"00CDA5",X"01BCA1",X"05B9A0",X"0FC1A7",X"0BBC9F",X"00BD99",X"12C6A9",X"2BBF9D",X"00513C",X"020109",X"1C0414",X"372032",X"5A2342",X"6D3454",X"612C46",X"040000",X"64390F",X"9F6639",X"3F190E",X"0B000B",X"0D2D42",X"2875A9",X"1F7EDC",X"0670E0",X"007CF0",X"007BEF",X"0877EA",X"0B74E7",X"207BE4",X"00307D",X"00022C",X"1C000D",X"530E2D",X"9D2660",X"C61C7D",X"D9078C",X"DC028D",X"D00F82",X"C11E77",X"7B235F",X"340414",X"0A0300",X"798322",X"ABAB25",X"807700",X"100900",X"030200",X"000600",X"09140C",X"293946",X"203759",X"314B7C",X"2C4A80",X"324F87",X"3F5D93",X"255070",X"234568",X"263D5F",X"2F3954",X"201F2F",X"130912",X"0A0005",X"0C000A",X"49323C",X"8D3B5F",X"AB1E63",X"D31E87",X"E3038A",X"F10085",X"FD098D",X"DF117D",X"981767",X"45001A",X"050308",X"060B11",X"0E0000",X"B65E3A",X"F5832B",X"F88109",X"FC720F",X"FE7600",X"FF7400",X"FC8527",X"B87035",X"0F0000",X"000409",X"7F8B77",X"F3FBF0",X"FAFDF4",X"FFFFFA",X"FFFFFA",X"FFFBFA",X"FDFBFE",X"FEFFFF",X"FAFDFF",X"F7FBFA",X"FFF7E1",X"DA964D",X"F1760C",X"FF7509",X"F57700",X"F57F03",X"F77611",X"FC8F10",X"D0713B",X"5F2001",X"140000",X"0A0300",X"8E7088",X"FFEBF4",X"EDFFFF",X"FFFAF4",X"FAFEFF",X"F4FEFF",X"FDFEFF",X"FFFBF9",X"FFFBFD",X"FBFEFF",X"ECF5FE",X"467CC4",X"0F6FBC",X"4179CC",X"264C7D",X"0E2D42",X"1E0F22",X"1F0000",X"883E0F",X"DF7931",X"E87522",X"D6790F",X"FFDDC7",X"FEFFFA",X"F6FFFF",X"FCFDF8",X"FFFDFE",X"FFFAFF",X"FFDBD4",X"CE9A68",X"96522D",X"080000",X"010002",X"617F59",X"80AF7B",X"74AE57",X"73AE52",X"90B361",X"5A6845",X"000005",X"765B54",X"FFE6D3",X"FDFEFF",X"FFFDFE",X"FFFEFF",X"FFFEFF",X"FEFEFE",X"FDFFFE",X"FFFFFF",X"FFFFFD",X"FEFDFB",X"F2FFFF",X"FBF3FE",X"F7FFFF",X"C8F3E9",X"3EAB8E",X"53908B",X"0D2A3A",X"00021B",X"082A81",X"256ED4",X"0B6BD9",X"0A6DD5",X"066AD9",X"0E68E0",X"0E5EC1",X"0E639C",X"C8EBE4",X"F1FFE6",X"FFF9FB",X"FFF6FF",X"FCFFF6",X"F8FFFF",X"FEFDFF",X"FFFBC1",X"F3E17D",X"A7A74F",X"000400",X"272123",X"200000",X"B06224",X"E68824",X"F3912C",X"E08F40",X"4D2F0B",X"190000",X"E3E4DE",X"FFFDF3",X"FBFFF2",X"F8FFFF",X"FFFCFF",X"F9FFFF",X"F5FBF7",X"FFFEF8",X"FFF8FB",X"F6F1F7",X"A27282",X"6F1940",X"71285D",X"571B37",X"37172F",X"0D0C2B",X"00012C",X"00003F",X"000F61",X"032F88",X"0D4AA5",X"1A5ABC",X"1169CD",X"0066D3",X"0166DA",X"0664D8",X"0565D5",X"1274DF",X"0F71DE",X"1F47A7",X"001241",X"0B0014",X"660F44",X"B61C7A",X"C50373",X"D90277",X"D70077",X"C90068",X"C9066C",X"AD1C69",X"35001D",X"000602",X"6A8F6D",X"75AF75",X"5CAA5F",X"5D9F55",X"67A35D",X"5F9351",X"6CA463",X"62A361",X"599F59",X"66A861",X"599450",X"669E61",X"649E4A",X"5F8949",X"020804",X"010007",X"90543C",X"E8863D",X"EA7E1B",X"FC8F2A",X"F07927",X"F68E47",X"975C30",X"0A0000",X"040700",X"91833C",X"D0A930",X"D3B51F",X"CFA805",X"D7AF0F",X"CAAB13",X"E0BA19",X"E4B716",X"C0A33D",X"222105",X"010700",X"58153E",X"C33088",X"CA0E6F",X"C40061",X"CA0171",X"CC097F",X"BF0776",X"C30E6B",X"9E0C5F",X"3F002B",X"211730",X"1B2E35",X"000518",X"000029",X"000035",X"00184B",X"000D44",X"000848",X"002570",X"093C8F",X"1454AE",X"175DBF",X"145DC3",X"215EBB",X"002471",X"000136",X"5A4C6D",X"3D1635",X"681A4C",X"9F1B6F",X"BE127E",X"CC046F",X"BE0974",X"C3117F",X"D00F7C",X"C70566",X"A01058",X"490A37",X"1B1732",X"00021B",X"C5DCEC"),
(X"FDFCF8",X"E8848E",X"D50000",X"E51836",X"CE011F",X"D50127",X"D90028",X"D70127",X"DD0028",X"D40229",X"DF0832",X"C2052D",X"3B1112",X"050001",X"0D3E38",X"2BB79A",X"13CBA5",X"00C8A0",X"05C0A5",X"01B59C",X"0BBDA3",X"0FC0A3",X"07CBA7",X"08BC9F",X"3BCFAD",X"31947F",X"0B0A12",X"0F0007",X"1D0618",X"25000D",X"300017",X"2B0010",X"090500",X"8C6137",X"DCA376",X"472116",X"0E020E",X"00091E",X"024F83",X"1978D6",X"0C76E6",X"0072E6",X"0079ED",X"006EE1",X"0C75E8",X"1B76DF",X"3C6DBA",X"1A2650",X"19000A",X"2D0007",X"67002A",X"C21879",X"D50388",X"DE048F",X"D41386",X"AA0760",X"711955",X"200000",X"615A2E",X"DAE483",X"FAFA74",X"E3DA57",X"BCB567",X"706F5D",X"414932",X"000500",X"000310",X"000729",X"000233",X"000F45",X"000C44",X"000339",X"000F2F",X"000629",X"000628",X"00001B",X"00000E",X"060005",X"150510",X"0B0009",X"321B25",X"722044",X"B12469",X"CB167F",X"E6068D",X"FF0095",X"F60286",X"D20470",X"A92878",X"85305A",X"020005",X"0B1016",X"0B0000",X"A14925",X"F6842C",X"F27B03",X"F86E0B",X"FF8309",X"FF830E",X"EB7416",X"B26A2F",X"342218",X"000409",X"97A38F",X"F7FFF4",X"FAFDF4",X"FFFFFA",X"FFFFFA",X"FFFDFC",X"FFFEFF",X"FBFCFF",X"FAFDFF",X"FCFFFF",X"D2C0AA",X"AD6920",X"FB8016",X"FF780C",X"F87A02",X"F98307",X"FC7B16",X"EE8102",X"E98A54",X"B27354",X"69503A",X"070000",X"E1C3DB",X"FFF8FF",X"EBFFFF",X"FFFBF5",X"FBFFFF",X"F5FFFF",X"FDFEFF",X"FFFBF9",X"FFFBFD",X"FBFEFF",X"ECF5FE",X"366CB4",X"004693",X"1850A3",X"00194A",X"000D22",X"08000C",X"73493D",X"C87E4F",X"E37D35",X"EA7724",X"D6790F",X"FFDCC6",X"FDFEF9",X"F6FFFF",X"FDFEF9",X"FFFDFE",X"FFF6FF",X"FFEEE7",X"E5B17F",X"5D1900",X"0E0402",X"09070A",X"6F8D67",X"7DAC78",X"6BA54E",X"72AD51",X"A0C371",X"4E5C39",X"000005",X"250A03",X"E8C7B4",X"FEFFFF",X"FFFCFD",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FFFFFF",X"FEFEFC",X"FFFEFC",X"E9FBFF",X"FFFBFF",X"F5FFFF",X"B3DED4",X"148164",X"00231E",X"000C1C",X"091932",X"385AB1",X"1E67CD",X"0363D1",X"0366CE",X"096DDC",X"1872EA",X"0757BA",X"58ADE6",X"DAFDF6",X"F8FFED",X"FFFBFD",X"FFF6FF",X"FCFFF6",X"F8FFFF",X"FFFEFF",X"FFFDC3",X"D8C662",X"414100",X"000400",X"040000",X"82593D",X"DC8E50",X"E0821E",X"FA9833",X"E89748",X"997B57",X"140000",X"E5E6E0",X"FFFCF2",X"FBFFF2",X"F7FEFF",X"FFFCFF",X"F6FCFF",X"F7FDF9",X"FFFCF6",X"FFFAFD",X"FFFAFF",X"865666",X"380009",X"4C0338",X"270007",X"17000F",X"0B0A29",X"101F4A",X"233575",X"334C9E",X"335FB8",X"2A67C2",X"1959BB",X"0860C4",X"016AD7",X"056ADE",X"0866DA",X"0A6ADA",X"0A6CD7",X"096BD8",X"375FBF",X"10305F",X"070010",X"520030",X"A60C6A",X"CC0A7A",X"D50073",X"D40074",X"D0026F",X"C8056B",X"AD1C69",X"4E1236",X"070D09",X"4D7250",X"649E64",X"49974C",X"60A258",X"69A55F",X"84B876",X"5B9352",X"6CAD6B",X"4E944E",X"64A65F",X"6EA965",X"679F62",X"619B47",X"729C5C",X"323834",X"010007",X"945840",X"E38138",X"F98D2A",X"DF720D",X"FF8836",X"E9813A",X"C88D61",X"433532",X"414439",X"6B5D16",X"CBA42B",X"D6B822",X"DCB512",X"D8B010",X"C6A70F",X"D2AC0B",X"DDB00F",X"C6A943",X"68674B",X"000300",X"45022B",X"BD2A82",X"D11576",X"CE056B",X"CF0676",X"C60379",X"BD0574",X"BF0A67",X"A81669",X"6E205A",X"332942",X"05181F",X"182033",X"080B34",X"18215A",X"143C6F",X"1B4077",X"2F5191",X"2C539E",X"2A5DB0",X"1858B2",X"1D63C5",X"165FC5",X"1754B1",X"3F66B3",X"364075",X"060019",X"27001F",X"4F0133",X"941064",X"B70B77",X"BE0061",X"BA0570",X"BF0D7B",X"CE0D7A",X"D91778",X"B2226A",X"672855",X"18142F",X"00021B",X"C6DDED"),
(X"FFF9FD",X"E68691",X"CF0000",X"E51934",X"D00020",X"D1032A",X"D20129",X"D30126",X"D70029",X"D00429",X"E30430",X"CE032E",X"5A0D15",X"070000",X"0E362D",X"46AC96",X"15C49D",X"00CD9F",X"07C9A7",X"00B79B",X"0ABEA1",X"08B599",X"06C1A2",X"07BEA2",X"00B299",X"1CD3B5",X"139885",X"004339",X"001710",X"000C0C",X"000A0B",X"10100E",X"0B0000",X"C2741F",X"F7971F",X"AD6510",X"501500",X"190001",X"010C2C",X"28456D",X"4179C4",X"267AD0",X"1372DC",X"026AE3",X"007AF6",X"0078F1",X"0E76E5",X"1475D6",X"003266",X"000835",X"040524",X"350D2F",X"8E255D",X"B9276E",X"8E275C",X"30172C",X"423C3E",X"312A00",X"D8CF34",X"F4EC1F",X"EFE507",X"F9EF11",X"FCED20",X"F6E12C",X"F4E54A",X"C1B71A",X"A7A10B",X"626200",X"131500",X"060800",X"010600",X"0D1100",X"07060C",X"1A0808",X"270000",X"8B4F1D",X"B16C21",X"B26E1B",X"874700",X"460A00",X"300000",X"1B0000",X"3C0C24",X"8A275E",X"CA2D7A",X"CF0D6D",X"E10C82",X"E6068D",X"CE1467",X"841245",X"010004",X"171516",X"080000",X"763A22",X"E37D33",X"FA7B06",X"F27908",X"FA8100",X"FF8105",X"F07C0D",X"CF7421",X"320300",X"000200",X"D5D1C6",X"FFFEFF",X"FBFBFD",X"FFFFFB",X"FDFDF5",X"FFFFF8",X"FFFFFD",X"F8F9FD",X"FEFEFF",X"FAF7FF",X"9B8B7E",X"7C471B",X"DD7D30",X"EC7000",X"FB7300",X"FF750B",X"FF7001",X"FF790A",X"F3760C",X"FF8624",X"D97B21",X"957F71",X"E6F1F5",X"FFFBFF",X"FFF8F6",X"FEFEF6",X"F8FFFF",X"F3FFFF",X"FEFFFF",X"FFFCFF",X"FEFBFF",X"FEFDFF",X"F7F1F1",X"3C353C",X"05090A",X"190200",X"200000",X"300000",X"AA5419",X"E77826",X"F36E05",X"FF7A0E",X"FF730B",X"DF7700",X"FFDDC4",X"F9FFF6",X"FAFFFF",X"FFFDF5",X"FFFCFA",X"FFFAF9",X"FFFDFF",X"E3D0CA",X"310900",X"050200",X"13250B",X"759E62",X"7AB45D",X"79AE54",X"7BB05E",X"90AB68",X"525740",X"040002",X"6B381B",X"E19F6D",X"FFF4E2",X"FFFCF9",X"FFFDFC",X"FFFFFD",X"FEFFFF",X"FEFFFF",X"FDFDFD",X"FDFBFC",X"FFFDFE",X"FFFCFF",X"F2FFFB",X"E8F2E9",X"76A092",X"1D3F49",X"000430",X"001263",X"0A5FB0",X"0069D2",X"0968E0",X"006ADA",X"0373D9",X"0064DC",X"177EFE",X"0755A8",X"C0D4EF",X"FBFFFF",X"FFFDFA",X"FFF5FF",X"FFF6FF",X"FDFEF6",X"F7FFFF",X"FDFDFF",X"FCF8DD",X"8A8164",X"000500",X"130C1C",X"5E1F00",X"DB7810",X"EB8614",X"EF870A",X"F97D09",X"FF8423",X"ED8A47",X"8A3A00",X"F8E9D2",X"FEFEF4",X"F7FFF8",X"F9FDFF",X"FFFDF9",X"FCFFFF",X"FDFEFF",X"FEFAF9",X"FEFFFA",X"F2FFFF",X"52617E",X"000033",X"002961",X"043695",X"0B4CAA",X"0F5FBE",X"0C62C5",X"0A61CA",X"0C64D0",X"0769D6",X"0069D6",X"0A5EDA",X"005DC1",X"0B6EC9",X"0A66D3",X"0258CF",X"0560CB",X"0163C8",X"0769D4",X"2369ED",X"1760AD",X"000D30",X"15092F",X"601357",X"B1167C",X"D30778",X"D2036F",X"C40169",X"D80671",X"C50767",X"841152",X"0D000B",X"395D4F",X"84B393",X"8DB68E",X"7D9B77",X"839E7D",X"6F8A6B",X"143113",X"779676",X"779C73",X"669062",X"6E9D69",X"6BA05A",X"699E5A",X"85AD6E",X"55814E",X"0E0300",X"0B0003",X"996244",X"EB8F42",X"FA7F31",X"F4891F",X"FF8E30",X"FA843C",X"9B5017",X"312316",X"000200",X"A19A63",X"C6B92C",X"CBB20D",X"C6A800",X"C9AC0A",X"CFA707",X"DBA908",X"CEAB2D",X"A5974C",X"001300",X"3A1B3A",X"841768",X"AC0766",X"C30569",X"D00578",X"CC007A",X"CA0076",X"BC0068",X"CE0975",X"C21D79",X"731A52",X"18001E",X"221F4E",X"143680",X"1560BD",X"1267C4",X"1969CC",X"155FC8",X"1360CC",X"0053C3",X"0965D4",X"0A68D9",X"0E6CDE",X"0A6EDD",X"0A6DCA",X"0F6AB1",X"24659B",X"000332",X"050025",X"250125",X"471936",X"A33F85",X"AB257C",X"AE046E",X"CB0A7D",X"D10072",X"C3005F",X"AE1661",X"721544",X"140000",X"CED9DD"),
(X"FFF8FC",X"E68691",X"CF0000",X"E51934",X"D10121",X"D2042B",X"D4032B",X"D50328",X"D70029",X"CF0328",X"DA0027",X"DA0F3A",X"5D1018",X"070000",X"001C13",X"2E947E",X"18C7A0",X"00C99B",X"01C3A1",X"09C0A4",X"09BDA0",X"01AE92",X"01BC9D",X"08BFA3",X"18D4BB",X"0DC4A6",X"41C6B3",X"47A49A",X"47928B",X"588080",X"364041",X"000000",X"372B13",X"E49641",X"F09018",X"E69E49",X"C98E6E",X"1F0007",X"000828",X"000931",X"013984",X"297DD3",X"1978E2",X"0870E9",X"0076F2",X"0074ED",X"0870DF",X"1273D4",X"296B9F",X"123360",X"020322",X"1F0019",X"590028",X"A21057",X"6E073C",X"170013",X"0A0406",X"867F37",X"EEE54A",X"EBE316",X"F4EA0C",X"F4EA0C",X"F3E417",X"FFEB36",X"E9DA3F",X"F2E84B",X"F4EE58",X"DEDE5C",X"C0C261",X"B8BA7B",X"B6BB93",X"5E6247",X"010006",X"0D0000",X"8A614D",X"CF9361",X"E19C51",X"E6A24F",X"D2924A",X"D19559",X"A37158",X"270200",X"210009",X"540028",X"A70A57",X"D51373",X"E10C82",X"DF0086",X"D71D70",X"7E0C3F",X"0B090E",X"0C0A0B",X"080000",X"571B03",X"D87228",X"FB7C07",X"F87F0E",X"FF8705",X"FC7A00",X"F27E0F",X"F39845",X"4D1E00",X"5C615D",X"FFFBF0",X"FFFEFF",X"FCFCFE",X"FFFFFB",X"FCFCF4",X"FFFFF8",X"FFFFFD",X"F8F9FD",X"FEFEFF",X"E3E0FD",X"190900",X"5A2500",X"DF7F32",X"FF8D19",X"FF7800",X"FE6B01",X"FF6700",X"FD7708",X"F77A10",X"FA7816",X"D3751B",X"EDD7C9",X"F4FFFF",X"FFF9FF",X"FFFCFA",X"FFFFF8",X"F8FFFF",X"F3FFFF",X"FEFFFF",X"FFFCFF",X"FEFBFF",X"FEFDFF",X"F7F1F1",X"342D34",X"000102",X"311A14",X"744B2F",X"AD7546",X"DC864B",X"E87927",X"FF7E15",X"FF7A0E",X"FF720A",X"DE7600",X"FFDCC3",X"F9FFF6",X"FAFFFF",X"FFFDF5",X"FFFCFA",X"FFF8F7",X"FFFBFD",X"FFF7F1",X"785046",X"0B0800",X"4E6046",X"80A96D",X"70AA53",X"73A84E",X"80B563",X"9BB673",X"464B34",X"070105",X"8E5B3E",X"C48250",X"FBE4D2",X"FFFEFB",X"FFFDFC",X"FFFFFD",X"FEFFFF",X"FEFFFF",X"FDFDFD",X"FDFBFC",X"FFFCFD",X"FFF8FD",X"EDFEF6",X"D9E3DA",X"042E20",X"00141E",X"24416D",X"3B50A1",X"156ABB",X"046DD6",X"0968E0",X"0F79E9",X"0061C7",X"0C70E8",X"005EDE",X"3E8CDF",X"E7FBFF",X"FAFEFF",X"FFFCF9",X"FFF3FF",X"FFF8FF",X"FEFFF7",X"F6FEFF",X"FCFCFF",X"FAF6DB",X"4A4124",X"000500",X"04000D",X"9B5C30",X"EF8C24",X"F38E1C",X"F99114",X"FD810D",X"F97312",X"EA8744",X"DF8F48",X"F6E7D0",X"FFFFF5",X"F8FFF9",X"F7FBFF",X"FFFEFA",X"FCFFFF",X"FBFCFF",X"FFFDFC",X"FFFFFB",X"EDFBFE",X"677693",X"1B2F62",X"2A538B",X"2E60BF",X"2566C4",X"1767C6",X"0F65C8",X"0E65CE",X"1068D4",X"0A6CD9",X"016BD8",X"0D61DD",X"005DC1",X"0568C3",X"0864D1",X"065CD3",X"0A65D0",X"0A6CD1",X"0D6FDA",X"1359DD",X"2E77C4",X"00284B",X"45395F",X"74276B",X"9C0167",X"D70B7C",X"D0016D",X"C5026A",X"D3016C",X"C70969",X"911E5F",X"220D20",X"25493B",X"88B797",X"91BA92",X"63815D",X"526D4C",X"163112",X"000F00",X"163515",X"759A71",X"739D6F",X"659460",X"6A9F59",X"689D59",X"85AD6E",X"6D9966",X"241915",X"080000",X"642D0F",X"D67A2D",X"FF8537",X"E4790F",X"FB8A2C",X"FA843C",X"BE733A",X"241609",X"121814",X"655E27",X"C5B82B",X"C2A904",X"CCAE00",X"C1A402",X"DAB212",X"C59300",X"D6B335",X"B4A65B",X"000B00",X"190019",X"B44798",X"BF1A79",X"C30569",X"C80070",X"C70075",X"D0037C",X"C1036D",X"CB0672",X"A90460",X"973E76",X"4B2D51",X"00002A",X"294B95",X"115CB9",X"075CB9",X"0F5FC2",X"0C56BF",X"1E6BD7",X"0B5FCF",X"1D79E8",X"0563D4",X"005DCF",X"0165D4",X"2689E6",X"025DA4",X"4D8EC4",X"284372",X"0A002A",X"341034",X"1D000C",X"8F2B71",X"C84299",X"B00670",X"C30275",X"DD087E",X"E71A83",X"B41C67",X"8D305F",X"1C0003",X"C6D1D5"),
(X"FFF9FF",X"E08992",X"C50500",X"DA1F34",X"CB0423",X"D4022F",X"D5022D",X"CF0628",X"D5072E",X"CE062B",X"DA0025",X"DA1237",X"8F0B20",X"320000",X"070000",X"154B3D",X"43B39B",X"0EBD96",X"01B393",X"0EC2A5",X"00BE9C",X"07BA9C",X"07C0A1",X"04BCA2",X"0ADBBE",X"03CAAD",X"04D0AD",X"1ECFB2",X"29D2B1",X"3DBC9F",X"325247",X"000700",X"9E561C",X"FD9027",X"FF8001",X"FC8F16",X"EF9D2F",X"955815",X"230000",X"1A0E00",X"0C091A",X"143E54",X"3179B4",X"1276D8",X"007AE2",X"0A78DA",X"0969DA",X"0070F4",X"136BE9",X"1C7CE0",X"004587",X"000532",X"1A042A",X"2B001B",X"311524",X"060006",X"001500",X"CBCE41",X"FFF017",X"FFDF00",X"FFDB01",X"FDE312",X"FFE70B",X"F5DA00",X"FFE500",X"FFE407",X"F8DE03",X"FFF911",X"FCF10C",X"FBF046",X"DBCA85",X"0F0007",X"17170F",X"0B0000",X"AA875D",X"E4AC59",X"E3971D",X"EC9000",X"F58C00",X"FF930B",X"F59C34",X"D7843E",X"6A3113",X"140000",X"2B0E13",X"651A3B",X"B0296E",X"C91D7F",X"CB3773",X"933B63",X"000200",X"0F0000",X"120800",X"0E0000",X"AA673A",X"F78127",X"F17103",X"FE8206",X"FD7200",X"F67300",X"FF8827",X"94370E",X"CBB3AF",X"FFF0F8",X"FEFCFF",X"FCFBFF",X"FFFFFF",X"FDFDFB",X"FDFDFB",X"FFFFFD",X"FBFDFA",X"FEFFFF",X"A0B1B9",X"000200",X"0D0000",X"7B5639",X"DB954F",X"DE6F15",X"FF7B18",X"FF7D00",X"F46F06",X"FF7602",X"FF7811",X"D3862C",X"F1E0C4",X"FFFFF4",X"FFFBFF",X"FDFEFF",X"FFFDFD",X"F9FFFF",X"F8FFFF",X"FFFEFB",X"FFFCFF",X"F9FDFF",X"FEFEFF",X"FFF0E0",X"AC631E",X"C5600E",X"DE7816",X"EA7C1A",X"FF8821",X"EA6C00",X"FF7900",X"FF7200",X"FF7900",X"FF6F08",X"DE7600",X"FFDFC2",X"F8FFF0",X"FBFFFF",X"FFFDF9",X"FFFEFA",X"FEFFF4",X"EAFFF7",X"FCFFFF",X"8A8D86",X"000B00",X"689A5F",X"80AF69",X"6AAC48",X"7DB25A",X"7DB470",X"829869",X"252317",X"251110",X"B26328",X"E37A1E",X"FDC18B",X"FFFEF8",X"FFFFFA",X"FFFEFC",X"FEFFFF",X"FEFFFF",X"FEFEFF",X"FEFCFF",X"FFFAFE",X"FDFFF4",X"FEFFFD",X"828894",X"000023",X"00245D",X"0156A9",X"0971E0",X"0864EB",X"006DD3",X"006FDB",X"0463D7",X"1971DF",X"1B81E6",X"064DA9",X"A1B3E5",X"FCFBF7",X"FFF8FF",X"FFF7FF",X"FFF7FF",X"FFFEFD",X"FEFFF9",X"FBFBFF",X"FFFCFF",X"F9F5EC",X"4B464C",X"100000",X"70321B",X"EC8025",X"FF8201",X"F17A02",X"EF7D03",X"FB7D19",X"ED790A",X"FF902D",X"F28C10",X"F6E4C0",X"F9FFFF",X"F9FFFF",X"F9F6FF",X"FFFFF1",X"FDFEF6",X"FDFAFF",X"FEFDFF",X"FEFFFA",X"F2F7FF",X"6583CC",X"124FB9",X"296DDC",X"0D6ED7",X"0766D2",X"0560D2",X"0661D6",X"0563D7",X"0464D5",X"0166D2",X"0368D0",X"086CE6",X"0363D3",X"005BC7",X"0263D4",X"0467DE",X"0768D9",X"0F6CD4",X"0760C8",X"1569BF",X"2E72BB",X"36578A",X"081535",X"0E0022",X"871C6A",X"C00C77",X"C2086D",X"D00B74",X"C30065",X"CD0E76",X"AF1D72",X"732F60",X"1F1E2C",X"4C635D",X"334036",X"151D20",X"001511",X"000E07",X"001710",X"000E08",X"556354",X"84AD8D",X"529768",X"5FA75B",X"588A55",X"589A5A",X"7FAD64",X"4D7946",X"000504",X"0C0800",X"A46843",X"E87838",X"E67E01",X"F27B03",X"FF7E29",X"FF9236",X"874B0C",X"3D241D",X"4B3C41",X"7E782C",X"BDAF34",X"C1AA0C",X"CEB10F",X"D1AB0C",X"CB9E00",X"D5AD1A",X"CFB137",X"433101",X"040000",X"655174",X"B963A4",X"AD0461",X"CF006C",X"D91382",X"AE0968",X"C80E71",X"C90064",X"CC096F",X"840B4E",X"361037",X"010F3C",X"1D4E9A",X"0C5ABF",X"0C6DD6",X"0461CB",X"065ECA",X"025DC6",X"0260C4",X"0D6ECC",X"0D6BC5",X"106AC2",X"257BE2",X"0558C0",X"075CC6",X"035CC2",X"3287E1",X"044388",X"00022E",X"040019",X"030010",X"5E425B",X"903E6E",X"AE2170",X"B20872",X"CD2594",X"C91882",X"DB167F",X"78002C",X"F6C0E0"),
(X"FFFAFF",X"E08992",X"C50500",X"DA1F34",X"CA0322",X"D3012E",X"D3002B",X"CD0426",X"D1032A",X"CD052A",X"DF002A",X"D0082D",X"A21E33",X"4E1319",X"080000",X"001709",X"1C8C74",X"25D4AD",X"0ABC9C",X"02B699",X"04C3A1",X"0EC1A3",X"00B495",X"0BC3A9",X"00C4A7",X"13DABD",X"04D0AD",X"0ABB9E",X"19C2A1",X"22A184",X"000F04",X"000600",X"BD753B",X"FE9128",X"FF8708",X"FA8D14",X"E89628",X"C38643",X"67432D",X"0A0000",X"0C091A",X"000B21",X"014984",X"197DDF",X"007AE2",X"0E7CDE",X"1070E1",X"0072F6",X"1971EF",X"0D6DD1",X"3081C3",X"2B4C79",X"0F001F",X"2E011E",X"150008",X"080108",X"ADC287",X"F3F669",X"F7DE05",X"FFE000",X"FFEA10",X"FBE110",X"F9E105",X"FFE601",X"FCE000",X"FFE70A",X"FDE308",X"F0DE00",X"F0E500",X"ECE137",X"796823",X"190111",X"14140C",X"150800",X"5A370D",X"C48C39",X"F6AA30",X"F99D0C",X"FC9303",X"FF8F07",X"E99028",X"ED9A54",X"B57C5E",X"391E15",X"140000",X"45001B",X"840042",X"BA0E70",X"BE2A66",X"7F274F",X"040700",X"7C695B",X"71675B",X"100000",X"7F3C0F",X"F27C22",X"FC7C0E",X"FC8004",X"FF7B06",X"FF810D",X"FA7A19",X"C76A41",X"F4DCD8",X"FFF4FC",X"FBF9FE",X"FDFCFF",X"FFFFFF",X"FFFFFD",X"FBFBF9",X"FEFEFC",X"FEFFFD",X"F5F7F6",X"71828A",X"020701",X"32241B",X"240000",X"A6601A",X"F8892F",X"FF7B18",X"F87100",X"F9740B",X"FF6F00",X"F66400",X"F8AB51",X"FFFADE",X"F9F5EA",X"FFFBFF",X"FBFCFF",X"FFFDFD",X"F9FFFF",X"F8FFFF",X"FFFEFB",X"FFFCFF",X"F9FDFF",X"FEFEFF",X"FFF0E0",X"DB924D",X"E6812F",X"E37D1B",X"ED7F1D",X"E76C05",X"F97B03",X"FF7E00",X"FF7800",X"FF7700",X"FF6F08",X"DE7600",X"FFE0C3",X"F9FFF1",X"FBFFFF",X"FFFDF9",X"FFFEFA",X"FEFFF4",X"EAFFF7",X"FCFFFF",X"D0D3CC",X"4C623B",X"8ABC81",X"79A862",X"6CAE4A",X"6FA44C",X"7DB470",X"748A5B",X"080600",X"0E0000",X"AD5E23",X"D56C10",X"F4B882",X"FFFCF6",X"FFFEF9",X"FFFEFC",X"FDFFFE",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFAFE",X"FFFFF6",X"E2E4E1",X"454B57",X"000025",X"245891",X"156ABD",X"0169D8",X"0460E7",X"0474DA",X"006FDB",X"0867DB",X"0F67D5",X"0C72D7",X"0B52AE",X"DBEDFF",X"FFFFFB",X"FFFAFF",X"FFF7FF",X"FFF8FF",X"FFFEFD",X"FAFBF5",X"F9F9FF",X"FFFDFF",X"F9F5EC",X"413C42",X"0E0000",X"AA6C55",X"F3872C",X"FD8000",X"FD860E",X"FC8A10",X"F27410",X"FF8E1F",X"F78522",X"E57F03",X"FEECC8",X"F9FFFF",X"F9FFFF",X"FDFAFF",X"FFFFF1",X"FCFDF5",X"FFFDFF",X"F9F8FD",X"FAFBF6",X"F7FCFF",X"6280C9",X"0D4AB4",X"2F73E2",X"0566CF",X"0463CF",X"0964D6",X"0E69DE",X"0A68DC",X"0464D5",X"0368D4",X"0A6FD7",X"0468E2",X"0C6CDC",X"005ECA",X"0061D2",X"0164DB",X"0061D2",X"0C69D1",X"0861C9",X"196DC3",X"185CA5",X"133467",X"041131",X"0E0022",X"6B004E",X"C5117C",X"C80E73",X"CC0770",X"CE0470",X"C6076F",X"AA186D",X"743061",X"1A1927",X"061D17",X"000500",X"000205",X"1D3A36",X"44716A",X"274C45",X"000802",X"000C00",X"6D9676",X"79BE8F",X"50984C",X"699B66",X"60A262",X"6D9B52",X"6D9966",X"0B1514",X"060200",X"783C17",X"EF7F3F",X"EF870A",X"F37C04",X"FF741F",X"FF9236",X"B67A3B",X"331A13",X"2D1E23",X"595307",X"CBBD42",X"C4AD0F",X"D0B311",X"CBA506",X"DFB211",X"CBA310",X"CFB137",X"867444",X"050100",X"402C4F",X"B05A9B",X"B30A67",X"DF0B7C",X"C70170",X"BD1877",X"C3096C",X"D4026F",X"CD0A70",X"9D2467",X"39133A",X"00002C",X"144591",X"1D6BD0",X"0869D2",X"0360CA",X"0961CD",X"0661CA",X"005EC2",X"096AC8",X"0260BA",X"0660B8",X"2076DD",X"1366CE",X"1065CF",X"1B74DA",X"176CC6",X"2362A7",X"2F4773",X"343049",X"090116",X"11000E",X"4F002D",X"9B0E5D",X"BD137D",X"B30B7A",X"B2016B",X"DE1982",X"8F1043",X"FBC5E5"),
(X"FFF8FF",X"E38593",X"C50300",X"D72034",X"CD0124",X"E10030",X"E1002D",X"D40227",X"D70028",X"D3022A",X"E3002B",X"CF0328",X"D50D34",X"9F102E",X"4E000E",X"000100",X"0E302F",X"40B69E",X"2DBFA8",X"08B599",X"02C8A4",X"07C0A0",X"00B192",X"0AC5AA",X"0BC8A8",X"04C8A4",X"0FC1A1",X"0ABF9C",X"30BAA0",X"3F5C5A",X"170000",X"664A3F",X"E6975C",X"E7A00A",X"FD9700",X"FF8100",X"EF8300",X"FF9F20",X"EE923D",X"935315",X"0D0000",X"2D2018",X"080007",X"1B2D53",X"3176C1",X"2676E9",X"0B65DD",X"007FDB",X"017AE5",X"0B70E6",X"0B6BE3",X"1581E4",X"0963AF",X"000F42",X"000823",X"00030C",X"827E59",X"D6D06E",X"EFE63F",X"EFE418",X"F0E809",X"EFEC00",X"FFF907",X"F2E400",X"EEE100",X"FDEE0D",X"FCEB17",X"EFDD23",X"FFF265",X"BCB05C",X"080100",X"130E12",X"3C0029",X"240017",X"230010",X"4C241C",X"B0834A",X"DB9C3F",X"E48F22",X"EC8617",X"FF9505",X"E48E03",X"F0A027",X"D27A23",X"520B00",X"1F0000",X"2A0809",X"3F0722",X"7B2F5D",X"360D2D",X"000A00",X"997658",X"736852",X"000908",X"290D00",X"CA703C",X"FF7A13",X"F37A09",X"F9760A",X"F07C05",X"ED790C",X"FFB57C",X"F5FFF1",X"F0FBFF",X"FCFBF9",X"FDFDFF",X"FCFBFF",X"FFFDFF",X"FBFBFF",X"FCFEFD",X"FEFFFA",X"DFE3D5",X"71A35C",X"2D4628",X"000500",X"040E0D",X"120003",X"B77457",X"F08C36",X"E97D0E",X"F57D0F",X"FF7F14",X"C76317",X"F7C5BE",X"FFF6EE",X"FFFAFE",X"F8FFFD",X"FCFFFF",X"FFFAFE",X"FFFEFF",X"FDFDFB",X"FFFDF6",X"FFFCFF",X"F6FEFF",X"FEFFFA",X"FFF0D1",X"F08A36",X"FE6100",X"FF7D05",X"FF780F",X"FE6E0E",X"FF8315",X"F77408",X"E86D0F",X"F77A02",X"FD7112",X"DD7802",X"FFE2C2",X"F8FFEA",X"FAFDFF",X"FFFDFF",X"F9FFFF",X"FFFAFF",X"F4FDF8",X"FFF6FF",X"E2F3EB",X"8AB077",X"6CB365",X"6DA05E",X"6EB660",X"88C069",X"82BC81",X"6B805F",X"040000",X"290E05",X"CE6E1A",X"F47200",X"F49F4E",X"F9F2EA",X"FFFBF5",X"FFFFFB",X"FDFFFE",X"FCFDFF",X"FFFEFF",X"FFFEFF",X"FFFBFF",X"F5F5FD",X"BEC5DF",X"000637",X"2065B0",X"2667CF",X"0968D4",X"006CD8",X"076BDB",X"0067D2",X"1270E4",X"126DDF",X"2E7DD9",X"193879",X"9794B3",X"FBFAFF",X"F2FFF8",X"FFFDFE",X"FCFBFF",X"F8FFF7",X"FAFFF3",X"F8F8FA",X"FDF6FF",X"FFFDFF",X"F4F2E6",X"2F2C1D",X"884808",X"FB882D",X"F7840F",X"F2810B",X"FD7C07",X"FA7900",X"FF8927",X"FF9616",X"E77E0B",X"ED8605",X"FFEFD8",X"FEFDFF",X"FEFFFD",X"FFFDFF",X"FEFEFC",X"FFFFF4",X"FFFBFF",X"F3FBFD",X"F8FFEC",X"F3FAFF",X"5181CB",X"0055BF",X"1C72DF",X"0D78D8",X"0669CF",X"025DCF",X"0461D8",X"086BE2",X"086BE0",X"0765D6",X"075DCE",X"0060C8",X"1366DC",X"1560D7",X"105FC4",X"1666BD",X"1E5CAF",X"274D96",X"2E477F",X"133950",X"1A1A50",X"210039",X"140019",X"130011",X"690040",X"C40473",X"CE0376",X"D4006D",X"D90A7C",X"C9006F",X"C6026E",X"A31164",X"480E37",X"00080D",X"0E3C2F",X"1C8A7F",X"29B49F",X"30C6AD",X"32988B",X"000C10",X"080002",X"485043",X"8AB997",X"70B370",X"5DA46A",X"6A975E",X"679C4C",X"6BA45D",X"436849",X"0B0000",X"472823",X"C9773F",X"F98424",X"FD7708",X"FA851C",X"EB8517",X"ED8820",X"B8672F",X"270000",X"5C5658",X"A49A5C",X"CEBB3A",X"BB9C03",X"D8B116",X"D3A80B",X"D5AA0D",X"D3A80E",X"DCA747",X"4B3400",X"070000",X"360E31",X"90306F",X"A51C6E",X"B31D74",X"AF1E6B",X"A91F6A",X"B52E7B",X"AA357C",X"7A2858",X"27001B",X"00011F",X"1A3B71",X"386BBC",X"1859AB",X"1A5AB1",X"1E5FBD",X"1D63C5",X"0B59BE",X"1D70D6",X"0A5BC4",X"0C59C1",X"0859C4",X"1A6DD3",X"075DC0",X"1C73DA",X"055AC5",X"0250B5",X"3A80D6",X"3275BC",X"00053F",X"151946",X"25153A",X"2A002D",X"791D6A",X"B72B8C",X"BB1675",X"C61A6E",X"A8005D",X"FFB6EB"),
(X"FFF7FF",X"E28492",X"C50300",X"D72034",X"CF0326",X"E30032",X"E40030",X"D7052A",X"D9002A",X"D8072F",X"E10029",X"D60A2F",X"CD052C",X"A91A38",X"560116",X"060805",X"000A09",X"0E846C",X"2CBEA7",X"19C6AA",X"00C29E",X"07C0A0",X"0EC9AA",X"00B89D",X"06C3A3",X"00BD99",X"11C3A3",X"10C5A2",X"159F85",X"000907",X"140000",X"5C4035",X"DA8B50",X"F0A913",X"F69000",X"FF8B08",X"FF930D",X"F39011",X"ED913C",X"D79759",X"706050",X"0A0000",X"180A17",X"000A30",X"003984",X"1E6EE1",X"1771E9",X"0085E1",X"017AE5",X"0C71E7",X"1070E8",X"0975D8",X"1F79C5",X"366194",X"12203B",X"00020B",X"080400",X"5D5700",X"ECE33C",X"FBF024",X"E8E001",X"F8F506",X"E7E100",X"FDEF06",X"F9EC08",X"F7E807",X"EBDA06",X"FFF036",X"E8D94C",X"625602",X"0A0300",X"1D181C",X"692556",X"6B305E",X"330220",X"200000",X"260000",X"9A5B00",X"F39E31",X"F48E1F",X"FA9000",X"F49E13",X"E99920",X"EA923B",X"D9925C",X"967156",X"180000",X"28000B",X"410023",X"360D2D",X"000A00",X"563315",X"443923",X"011110",X"160000",X"A94F1B",X"FF7C15",X"F57C0B",X"FE7B0F",X"F5810A",X"F37F12",X"FFC188",X"F1FEED",X"F7FFFF",X"FEFDFB",X"FEFEFF",X"F9F8FE",X"FFFDFF",X"FDFDFF",X"FDFFFE",X"FEFFFA",X"CED2C4",X"689A53",X"768F71",X"0C190F",X"000807",X"0E0000",X"480500",X"D6721C",X"F68A1B",X"F1790B",X"F36C01",X"F89448",X"FFE1DA",X"FFF8F0",X"FFFDFF",X"F0FBF5",X"FCFFFF",X"FFFAFE",X"FFFEFF",X"FDFDFB",X"FFFDF6",X"FFFCFF",X"F6FEFF",X"FEFFFA",X"FFF0D1",X"EE8834",X"FF6C0B",X"FB7300",X"FF7910",X"FF7313",X"F27204",X"F57206",X"F27719",X"F97C04",X"FF7314",X"DF7A04",X"FFE3C3",X"F7FFE9",X"F9FCFF",X"FFFDFF",X"F9FFFF",X"FFF6FF",X"F9FFFD",X"FFF9FF",X"F1FFFA",X"ACD299",X"5CA355",X"71A462",X"67AF59",X"87BF68",X"6EA86D",X"1D3211",X"040000",X"492E25",X"D47420",X"F87600",X"D07B2A",X"F1EAE2",X"FDF8F2",X"FFFFFB",X"FEFFFF",X"FCFDFF",X"FFFEFF",X"FFFEFF",X"FFFBFF",X"F5F5FD",X"8188A2",X"264E7F",X"2C71BC",X"1E5FC7",X"0564D0",X"0473DF",X"0A6EDE",X"0574DF",X"0A68DC",X"0560D2",X"1E6DC9",X"001051",X"CECBEA",X"F6F5FA",X"F4FFFA",X"FFFCFD",X"FBFAFF",X"F9FFF8",X"FBFFF4",X"FBFBFD",X"FFFAFF",X"FFFDFF",X"F1EFE3",X"6A6758",X"C38343",X"F68328",X"F5820D",X"F1800A",X"FF820D",X"FE7D00",X"FF8A28",X"EB8202",X"FD9421",X"E27B00",X"FFE9D2",X"FAF9FF",X"FEFFFD",X"FBF8FF",X"FFFFFD",X"FFFFF4",X"FBF3FF",X"F9FFFF",X"FBFFEF",X"EAF1FB",X"5181CB",X"015EC8",X"0C62CF",X"0772D2",X"086BD1",X"0661D3",X"025FD6",X"0164DB",X"0568DD",X"0967D8",X"0D63D4",X"0164CC",X"1164DA",X"1762D9",X"0C5BC0",X"1666BD",X"1553A6",X"001A63",X"000139",X"000A21",X"000036",X"2C0244",X"3D1A42",X"40223E",X"85185C",X"C0006F",X"CC0174",X"DC0175",X"CD0070",X"D30979",X"D20E7A",X"CC3A8D",X"420831",X"000409",X"427063",X"36A499",X"28B39E",X"1BB198",X"2E9487",X"3E5A5E",X"0B0005",X"000500",X"7DAC8A",X"7CBF7C",X"73BA80",X"77A46B",X"5F9444",X"70A962",X"5B8061",X"160606",X"160000",X"A6541C",X"FC8727",X"FF790A",X"F68118",X"E57F11",X"EE8921",X"E08F57",X"72433D",X"2A2426",X"574D0F",X"B5A221",X"D0B118",X"D7B015",X"DBB013",X"D2A70A",X"CA9F05",X"E0AB4B",X"8A733F",X"070000",X"31092C",X"6D0D4C",X"A01769",X"8C004D",X"890045",X"880049",X"8F0855",X"88135A",X"5B0939",X"27001B",X"0E0F2D",X"103167",X"1F52A3",X"0C4D9F",X"1454AB",X"2E6FCD",X"185EC0",X"1260C5",X"1669CF",X"1566CF",X"1360C8",X"1869D4",X"0052B8",X"1C72D5",X"055CC3",X"1166D1",X"0F5DC2",X"0B51A7",X"2265AC",X"465993",X"171B48",X"201035",X"491B4C",X"650956",X"A71B7C",X"C82382",X"C2166A",X"AA005F",X"FFB8ED"),
(X"FFFBFF",X"E28484",X"BB0700",X"EF1837",X"D10220",X"DA0B25",X"D50024",X"DC0039",X"DB002B",X"D4062D",X"CB0226",X"D40024",X"E5002D",X"DC0B35",X"99051D",X"530000",X"1B0102",X"070000",X"406860",X"4DB4A1",X"26B99F",X"1BBFA4",X"0FC3A6",X"0BD1AE",X"09BD9A",X"02C1A0",X"05B79D",X"35B2A0",X"226254",X"000D00",X"061208",X"000100",X"584211",X"CA964A",X"F79D2D",X"F68608",X"FE8C10",X"F78D15",X"F69012",X"F8940B",X"F39939",X"B36A26",X"280000",X"110000",X"000005",X"13324F",X"2B6CAE",X"227CDC",X"107AEA",X"0276DD",X"007AE1",X"0076E8",X"0068E7",X"1770E4",X"3076CC",X"003771",X"000631",X"06071B",X"62543A",X"E1CC79",X"FEED61",X"EBDD22",X"F9EC12",X"F3E601",X"EEEA05",X"F0E416",X"FFEE4D",X"C6B34D",X"414312",X"000100",X"23000E",X"7A003D",X"D1167F",X"DF1480",X"BC0D6C",X"640031",X"370015",X"160000",X"624A24",X"D79F6E",X"E69F33",X"EF9824",X"FE9013",X"FE8705",X"FF9F26",X"E78E2A",X"A46015",X"592200",X"180000",X"070002",X"0C0D12",X"040313",X"000023",X"000918",X"080700",X"563226",X"DF7B2D",X"F78018",X"F77300",X"F57D05",X"E08F3D",X"FFDECD",X"FFF8FF",X"FAFEFF",X"FCFFFF",X"FEFAF9",X"FFF9FF",X"FCFDFF",X"FBF9FC",X"FFFCF7",X"F1FDE5",X"8AB878",X"6DA76C",X"6FA35B",X"6E9552",X"000B00",X"070908",X"110001",X"563117",X"BE8D52",X"F77E2D",X"CD6E2A",X"ECB785",X"FFFDE1",X"F3F9EF",X"F7FFFF",X"FCFFFF",X"FFFBFF",X"FFFEFF",X"FFFFFD",X"FEFEFC",X"FEFFFD",X"FDFDFD",X"FFFBFA",X"FFFDF7",X"FAF4E8",X"FE852A",X"F27410",X"F36F00",X"FF7805",X"FF7502",X"FB6D01",X"FE730C",X"FE7610",X"FA7E02",X"FF7400",X"E47519",X"FFE4B1",X"F1FFF4",X"F8FFFF",X"FFFDFD",X"FBFEF5",X"F8FFED",X"FFFCFF",X"FFF7FF",X"F8F9F1",X"B8D9A2",X"6EA853",X"68A24E",X"8BBA74",X"82BB6A",X"90B07F",X"1D2B1E",X"040000",X"6A300B",X"EF7826",X"F9760E",X"DE750C",X"FFD9C3",X"FFFFE7",X"FFFCF9",X"FFF4FF",X"F7FFFF",X"FBFFFF",X"FFF4F9",X"FBFFFD",X"C8F4FF",X"1D5AB7",X"1C7AEE",X"006CCF",X"0068CF",X"026ED3",X"086FD4",X"096DE7",X"016DD9",X"1565C8",X"3863B1",X"081F4B",X"52626F",X"E9F3F2",X"FFFEFF",X"FFF7FF",X"FCFDFF",X"FFFFFF",X"FEFDF8",X"FEFFF5",X"FDFEFF",X"FFFCFF",X"FFFDFA",X"FCF3D2",X"D58F53",X"EB780D",X"FF921B",X"FF8D11",X"F97400",X"FE8012",X"F07800",X"F18D11",X"FF8C0E",X"F78E3D",X"BA6431",X"E1E0DC",X"FEFFFA",X"FFF7F0",X"FFFDFA",X"EFFFFF",X"F7FFFF",X"F6FDF6",X"FFFDFF",X"FFF6FA",X"EFFDFF",X"588CC8",X"0050C3",X"1069DD",X"0065E0",X"0D72E4",X"0061C7",X"0868CC",X"0664C8",X"0B61C4",X"1A65C2",X"1D5FB5",X"1B60A3",X"3961A7",X"3C4A89",X"262C5C",X"101938",X"07001F",X"1F001E",X"4C0038",X"7E0044",X"95115D",X"A1156E",X"AC1177",X"BB1080",X"C2077C",X"C70077",X"D7077F",X"CD0076",X"D10078",X"E20C88",X"CB0073",X"C61C7F",X"761353",X"06000E",X"366960",X"279F95",X"06A68C",X"00BB93",X"06AE8D",X"359E90",X"184644",X"000B07",X"404C40",X"65A372",X"5FA068",X"76B974",X"619F52",X"65994F",X"759A64",X"26381E",X"000300",X"623919",X"DA7A48",X"FB7629",X"F57A13",X"EC770E",X"FF8B30",X"FF853A",X"C35E1A",X"130000",X"21230B",X"757E49",X"C4B33F",X"C7A200",X"D7B013",X"C2A30B",X"D6B906",X"D7A11A",X"B18944",X"110300",X"030A1A",X"0E0210",X"3D0F1A",X"230000",X"0B0000",X"110000",X"0E0000",X"0E0100",X"0A0000",X"2B1F21",X"312732",X"07000F",X"120E1F",X"080E0E",X"020C16",X"202E48",X"203054",X"0E1D44",X"0C2043",X"213A63",X"294479",X"325994",X"315B95",X"2F5D98",X"2C5595",X"274991",X"2B4C93",X"38619F",X"1D5085",X"3D65AD",X"396099",X"162F57",X"1D203F",X"080019",X"340B35",X"A24C8B",X"B73387",X"761248",X"FFC0EA"),
(X"FFFAFF",X"DF8181",X"BB0700",X"EC1534",X"D0011F",X"D70822",X"D90128",X"DB0038",X"D80028",X"D2042B",X"CE0529",X"D80028",X"E4002C",X"D80731",X"A8142C",X"791A22",X"341A1B",X"060000",X"00140C",X"005643",X"11A48A",X"26CAAF",X"0EC2A5",X"0BD1AE",X"0FC3A0",X"12D1B0",X"14C6AC",X"1C9987",X"003729",X"001709",X"313D33",X"030500",X"150000",X"875307",X"F09626",X"FC8C0E",X"FB890D",X"FF9921",X"ED8709",X"FB970E",X"F19737",X"E39A56",X"8E623F",X"281205",X"101116",X"000E2B",X"003779",X"227CDC",X"0C76E6",X"0071D8",X"0072D9",X"007AEC",X"0572F1",X"166FE3",X"286EC4",X"3772AC",X"23325D",X"1A1B2F",X"150700",X"644F00",X"CEBD31",X"FFF53A",X"EEE107",X"FAED08",X"F0EC07",X"EDE113",X"F0DA39",X"513E00",X"040600",X"1C1D18",X"3A0225",X"A22665",X"D0157E",X"DA0F7B",X"C41574",X"A12A6E",X"581236",X"1D0000",X"1D0500",X"5C2400",X"CF881C",X"F29B27",X"FF9316",X"FF8F0D",X"FF9219",X"E68D29",X"E8A459",X"BF8850",X"2F1305",X"2B2026",X"000106",X"323141",X"43476D",X"132332",X"050400",X"210000",X"CC681A",X"F17A12",X"FF8000",X"ED7500",X"FFB361",X"FFF1E0",X"FFF3FF",X"FCFFFF",X"F3F7FA",X"FFFEFD",X"FFFBFF",X"F8F9FF",X"F5F3F6",X"FFFDF8",X"E1EDD5",X"81AF6F",X"6EA86D",X"7AAE66",X"7DA461",X"6A805A",X"1E201F",X"0E0000",X"1D0000",X"7F4E13",X"F07726",X"E48541",X"FFD5A3",X"FFFDE1",X"F9FFF5",X"F4FFFF",X"F9FCFF",X"FFFDFF",X"FFFEFF",X"FFFFFD",X"FEFEFC",X"FEFFFD",X"FDFDFD",X"FFFBFA",X"FFFDF7",X"FAF4E8",X"F67D22",X"F87A16",X"FD790A",X"FF7502",X"FE7100",X"FF770B",X"FF7B14",X"F8700A",X"F77B00",X"FF7C08",X"D7680C",X"FFE8B5",X"F5FFF8",X"F8FFFF",X"FDF7F7",X"FEFFF8",X"FCFFF1",X"FFF8FF",X"FFF5FF",X"FFFFF8",X"CBECB5",X"6AA44F",X"78B25E",X"76A55F",X"89C271",X"6D8D5C",X"000A00",X"040000",X"8E542F",X"F07927",X"FF7D15",X"D97007",X"FFD2BC",X"FFFFE8",X"FFFDFA",X"FFF6FF",X"F9FFFF",X"FBFFFF",X"FFF7FC",X"FBFFFD",X"A7D3EC",X"2663C0",X"0361D5",X"006ED1",X"0A7EE5",X"006ACF",X"0067CC",X"0063DD",X"006BD7",X"1969CC",X"305BA9",X"00022E",X"97A7B4",X"F8FFFF",X"F6F4F7",X"FFFAFF",X"FCFDFF",X"FFFFFF",X"FEFDF8",X"FEFFF5",X"FDFEFF",X"FFFBFF",X"FFFDFA",X"FBF2D1",X"DC965A",X"EE7B10",X"FB8E17",X"F48206",X"FF7F06",X"FC7E10",X"FD850D",X"E78307",X"FF8C0E",X"E9802F",X"5D0700",X"E7E6E2",X"FEFFFA",X"FFF7F0",X"FFFCF9",X"F1FFFF",X"F8FFFF",X"F7FEF7",X"FFFDFF",X"FFF5F9",X"EFFDFF",X"588CC8",X"0858CB",X"136CE0",X"0971EC",X"0D72E4",X"0B6ED4",X"0262C6",X"0E6CD0",X"0E64C7",X"1560BD",X"1052A8",X"094E91",X"072F75",X"000948",X"00002C",X"000322",X"1B1433",X"4D1B4C",X"761C62",X"9B1C61",X"A4206C",X"A71B74",X"AE1379",X"BB1080",X"C2077C",X"C50075",X"CE0076",X"D80B81",X"F12098",X"D00076",X"C5006D",X"BE1477",X"8D2A6A",X"100418",X"10433A",X"1F978D",X"05A58B",X"00B189",X"05AD8C",X"349D8F",X"43716F",X"000602",X"000500",X"498756",X"60A169",X"66A964",X"68A659",X"5B8F45",X"799E68",X"5B6D53",X"000300",X"290000",X"CF6F3D",X"FF7A2D",X"FF8A23",X"E77209",X"F8781D",X"F97F34",X"DD7834",X"503B28",X"010300",X"4F5823",X"B3A22E",X"D9B40E",X"CAA306",X"C6A70F",X"CDB000",X"EBB52E",X"AC843F",X"1A0C09",X"0F1626",X"403442",X"481A25",X"3F1517",X"45372C",X"4C382D",X"271606",X"423524",X"392C23",X"090000",X"060007",X"090011",X"01000E",X"020808",X"00020C",X"000D27",X"000125",X"05143B",X"000427",X"000D36",X"00073C",X"072E69",X"07316B",X"002661",X"022B6B",X"001058",X"03246B",X"07306E",X"05386D",X"113981",X"254C85",X"385179",X"191C3B",X"110022",X"260027",X"731D5C",X"AC287C",X"5E0030",X"FEBDE7"),
(X"F8FCFB",X"BC869D",X"88100F",X"CF203F",X"C90326",X"D20236",X"DE0230",X"DF0013",X"E0002D",X"DD002D",X"D8012B",X"D5022B",X"D0012B",X"CB022C",X"CB0832",X"CC0F39",X"89001A",X"5A0006",X"240000",X"000203",X"112929",X"4D6C6E",X"5F9E96",X"4AB19C",X"46C49E",X"1CBC98",X"3ED0BB",X"488C8D",X"000106",X"040800",X"84A37A",X"699361",X"000305",X"090601",X"725337",X"DA9C53",X"E99018",X"F98F00",X"FF9306",X"FB8B0D",X"FDA216",X"F59910",X"FCA82E",X"C27E2D",X"270000",X"0B0005",X"030923",X"1F3149",X"3575BF",X"2D74D0",X"1B6DDD",X"1070E9",X"056FE9",X"0370E7",X"0A76F2",X"016AEA",X"207AF4",X"0D53A9",X"002852",X"000712",X"000600",X"979C66",X"E7DB6F",X"F8DE49",X"F6D72E",X"FBEA78",X"757748",X"000300",X"2F1423",X"4A0015",X"B60F61",X"E00D82",X"E60078",X"E0067E",X"E0007D",X"E80787",X"B8006D",X"A41A67",X"630F33",X"160000",X"220006",X"98725D",X"CD9A5B",X"E8A43F",X"EA9619",X"FA9C18",X"FFA121",X"F4961C",X"D57C3A",X"7A4D30",X"000408",X"1D5087",X"2D75D9",X"0A4E9F",X"000927",X"0D0005",X"81432A",X"E27C3C",X"FF7C21",X"DA7003",X"FCCAB1",X"FEFEFF",X"EFFCF3",X"FFFDF0",X"FFFEFF",X"F8F8F6",X"FEF9FD",X"FFFDFF",X"FEFFF4",X"ECFFEC",X"ADD2A7",X"85B65B",X"7EAF5E",X"71AC58",X"6FB262",X"7FB373",X"6D8760",X"020600",X"090400",X"050100",X"582D0A",X"A8896D",X"FEEDDD",X"FFFDFA",X"FCFFFF",X"FAFFFF",X"F6F8F7",X"FFFFFA",X"FFFEFF",X"FFFFFD",X"FEFEFC",X"FFFFFF",X"FDFDFF",X"FFFBFA",X"FFFDF7",X"FAF4E8",X"FE7B23",X"F97310",X"FD7306",X"FF7400",X"FF6F00",X"FF7400",X"FF7C06",X"FE7902",X"F27A19",X"FC7E27",X"D27236",X"FEDAC0",X"FEFFFF",X"FAFDFF",X"FFFDFF",X"F5F7FF",X"FFFBFF",X"FEFFFF",X"F7F8FD",X"FDFDFF",X"F3FFED",X"7EA65D",X"73AA45",X"8CBD61",X"96AA65",X"55654A",X"000202",X"1C0000",X"C36D30",X"F97312",X"FF7C0D",X"E66E00",X"F7BF9A",X"FCFFF1",X"F9FFFF",X"FFFCFF",X"F7FFFF",X"FBFFFF",X"FFFCF9",X"EBFCFF",X"5FA9E6",X"1058C7",X"1565E2",X"0C68D7",X"0465DA",X"0366DB",X"0469D5",X"0869DE",X"1D63D2",X"365CA3",X"0A0F2C",X"060004",X"F0E6E7",X"FFFDFB",X"FFFFFA",X"F8FFFB",X"FDFFFE",X"FFFFFF",X"FEFDF9",X"FEFFF9",X"FCFDFF",X"FFFBFF",X"FFFDF7",X"FAF2CE",X"DD873C",X"FF8A26",X"F87F24",X"FE831B",X"F78100",X"F49310",X"F08618",X"F78235",X"B17A5C",X"4A3B28",X"130600",X"DEEBFE",X"FEF6FF",X"FFFEFA",X"F2F3ED",X"FFFFFF",X"FEFFFA",X"FAFFF8",X"FFFCFF",X"FFFAFF",X"EAFDFF",X"4F89C8",X"0757CA",X"0D62D9",X"106BD6",X"1963C4",X"2C64B7",X"285A9F",X"33649C",X"2D4F7D",X"1B2048",X"0E001F",X"130017",X"1A0018",X"370029",X"60003C",X"86004E",X"AE0965",X"CA0F76",X"CF0978",X"DA0174",X"D20274",X"C80175",X"C20375",X"C30778",X"C9097A",X"CF0978",X"D40A78",X"DA0B73",X"CE0B71",X"BF096D",X"C71978",X"BD2476",X"8B225A",X"310B24",X"081617",X"1F8A80",X"23AD96",X"04A788",X"00A686",X"01AB8E",X"23B398",X"044A40",X"0C070E",X"567162",X"93BA9D",X"5D9362",X"61A25E",X"63A158",X"679759",X"648058",X"031200",X"060004",X"8F6149",X"DD8848",X"FF9239",X"F77F0E",X"FA7F00",X"F37C06",X"EF8122",X"B85B1E",X"3D1516",X"423D3A",X"857132",X"D7B643",X"CBB71A",X"C6AF00",X"CB9B00",X"CAC10E",X"B5AE15",X"404000",X"050400",X"463548",X"AB7C6A",X"C4783A",X"D17427",X"E78440",X"F08342",X"E47138",X"C75F2C",X"D07E4C",X"C27B45",X"B05F28",X"B95C21",X"C56340",X"AF5533",X"A65B3C",X"7B4634",X"422426",X"1D1220",X"151918",X"000800",X"001000",X"16260B",X"2E3D20",X"010B00",X"020500",X"030100",X"0F0C00",X"040200",X"000C00",X"00100D",X"000F12",X"19262C",X"000D0E",X"334132",X"2A2B1D",X"43313F",X"1C000D",X"D5C5D2"),
(X"F9FDFC",X"B88299",X"7A0201",X"D32443",X"C90326",X"D10135",X"DD012F",X"E00114",X"E30030",X"DC002C",X"D60029",X"D4012A",X"D1022C",X"CA012B",X"C6032D",X"C60933",X"AC1C3D",X"92263E",X"481923",X"040809",X"000707",X"000B0D",X"002F27",X"005F4A",X"02805A",X"1BBB97",X"3BCDB8",X"206465",X"000005",X"6B6F60",X"97B68D",X"9DC795",X"3E494B",X"030000",X"190000",X"8E5007",X"EC931B",X"FE9404",X"FE8F02",X"FF981A",X"F4990D",X"F1950C",X"F09C22",X"E09C4B",X"B18369",X"200E1A",X"00001A",X"000B23",X"00317B",X"2168C4",X"2476E6",X"0969E2",X"127CF6",X"0976ED",X"0D79F5",X"0871F1",X"156FE9",X"2D73C9",X"406B95",X"2B4651",X"000600",X"050A00",X"504400",X"E2C833",X"FDDE35",X"968513",X"040600",X"0C130C",X"17000B",X"852650",X"BD1668",X"DE0B80",X"F70F89",X"DA0078",X"E0007D",X"E60585",X"D11786",X"B22875",X"782448",X"230B0B",X"1A0000",X"290300",X"723F00",X"BF7B16",X"E89417",X"F39511",X"F79818",X"FA9C22",X"F39A58",X"794C2F",X"000307",X"1F5289",X"2C74D8",X"2B6FC0",X"0A2745",X"100008",X"4C0E00",X"DD7737",X"FA751A",X"EE8417",X"FFD7BE",X"FEFEFF",X"F7FFFB",X"FFFEF1",X"FDFCFF",X"FFFFFD",X"FCF7FB",X"FFFDFF",X"F9FDEF",X"EEFFEE",X"9DC297",X"74A54A",X"84B564",X"72AD59",X"72B565",X"75A969",X"8EA881",X"898D7C",X"201B17",X"292522",X"260000",X"BFA084",X"FFFCEC",X"FCF8F5",X"F8FCFF",X"FAFFFF",X"FBFDFC",X"FFFFFA",X"FFFEFF",X"FFFFFD",X"FEFEFC",X"FFFFFF",X"FDFDFF",X"FFFBFA",X"FFFDF7",X"FAF4E8",X"FF7C24",X"F46E0B",X"FE7407",X"FF7A06",X"FF7300",X"FD7000",X"F77000",X"F67100",X"FB8322",X"EE7019",X"DA7A3E",X"FFEAD0",X"F9FBFA",X"F9FCFF",X"F9F6FF",X"FCFEFF",X"FFFDFF",X"F9FBFA",X"FEFFFF",X"FEFEFF",X"EBFAE5",X"9DC57C",X"74AB46",X"73A448",X"8CA05B",X"061600",X"040A0A",X"4F3222",X"C56F32",X"FD7716",X"FA7001",X"EF7706",X"E1A984",X"F8FCED",X"F9FFFF",X"FFFAFF",X"F6FFFF",X"F8FEFC",X"FFFEFB",X"DDEEFE",X"357FBC",X"0E56C5",X"1C6CE9",X"136FDE",X"0263D8",X"086BE0",X"0368D4",X"0263D8",X"1C62D1",X"02286F",X"00011E",X"6A6068",X"F7EDEE",X"FEF6F4",X"FFFFFA",X"EBF6EE",X"FEFFFF",X"FFFFFF",X"FFFEFA",X"FFFFFA",X"FCFDFF",X"FFFBFF",X"FFFDF7",X"FAF2CE",X"E58F44",X"FA7C18",X"F87F24",X"FB8018",X"FD8703",X"EB8A07",X"EF8517",X"E87326",X"551E00",X"0E0000",X"0B0000",X"D9E6F9",X"FFF9FF",X"FDF8F4",X"FFFFFA",X"FCFCFC",X"FDFEF9",X"FBFFF9",X"FEFBFF",X"FFFBFF",X"EAFDFF",X"4E88C7",X"0C5CCF",X"1065DC",X"0C67D2",X"1F69CA",X"1E56A9",X"0C3E83",X"001C54",X"000D3B",X"000026",X"160227",X"220726",X"40163E",X"6D285F",X"932D6F",X"A92271",X"B8136F",X"C60B72",X"CC0675",X"D2006C",X"CD006F",X"CB0478",X"C8097B",X"C30778",X"C50576",X"CC0675",X"CF0573",X"DA0B73",X"C10064",X"CD177B",X"BD0F6E",X"B01769",X"811850",X"350F28",X"000506",X"00695F",X"1CA68F",X"07AA8B",X"04AF8F",X"11BB9E",X"1CAC91",X"286E64",X"030005",X"000A00",X"638A6D",X"6EA473",X"5C9D59",X"619F56",X"6E9E60",X"85A179",X"4A5944",X"090007",X"582A12",X"D37E3E",X"EE8027",X"F67E0D",X"FF8A09",X"FC850F",X"F28425",X"D87B3E",X"694142",X"5A5552",X"4B3700",X"BA9926",X"D4C023",X"BAA300",X"DFAF0D",X"B3AA00",X"C2BB22",X"868630",X"010000",X"0A000C",X"A87967",X"E39759",X"E78A3D",X"E88541",X"F78A49",X"EE7B42",X"DD7542",X"EF9D6B",X"E59E68",X"DC8B54",X"DA7D42",X"DB7956",X"DD8361",X"EBA081",X"C5907E",X"4A2C2E",X"060009",X"1B1F1E",X"2D3A20",X"293B21",X"3D4D32",X"324124",X"0E1800",X"1C1F0E",X"514F42",X"524F3C",X"403E27",X"0C1D0D",X"000D0A",X"00070A",X"000309",X"000405",X"000600",X"27281A",X"342230",X"472438",X"E5D5E2"),
(X"FFF8FF",X"939194",X"380A00",X"C52A52",X"D60029",X"D50424",X"C90628",X"D40636",X"D1042F",X"D2012B",X"D4002B",X"D2032D",X"CF082F",X"CE0730",X"D3012E",X"D8002E",X"C70028",X"DA133E",X"B50B30",X"6D0010",X"380000",X"280000",X"220000",X"150000",X"0D0000",X"2B4C45",X"345C5B",X"000004",X"060700",X"568C52",X"73C271",X"7EBD6C",X"7DBC85",X"124620",X"000C00",X"080400",X"82593D",X"E09752",X"ED921D",X"F49200",X"FF8900",X"FE9005",X"FF9A1A",X"F89017",X"FF9D2F",X"CD721F",X"460B00",X"1B0000",X"060000",X"0F1835",X"4269AE",X"3079D5",X"0C70CE",X"0476D9",X"006FE2",X"0677FB",X"0082DA",X"007ADC",X"097EE7",X"237DDD",X"134E94",X"00143A",X"00030C",X"2B312D",X"686651",X"060100",X"090000",X"200011",X"8B195F",X"D50F7E",X"F80F84",X"E2016B",X"E60078",X"D30778",X"DE1484",X"DD0078",X"EB0484",X"EA0584",X"D2117E",X"91075D",X"390B16",X"0B0002",X"000909",X"000700",X"6A6547",X"AB8449",X"E0A046",X"E19827",X"F39756",X"A16D48",X"000004",X"1C4D87",X"2573E0",X"2577DD",X"265897",X"000533",X"080000",X"875323",X"C87412",X"F0A57B",X"FFF2D0",X"EEFFFF",X"F4FFFF",X"FFFAEA",X"FFFCFF",X"F6FBF4",X"FEFDF9",X"FFF4F3",X"FFFFF4",X"D6F7E6",X"7DAB87",X"86AF63",X"7CBA4F",X"79AF4F",X"7DAF58",X"83BE64",X"6DB051",X"74B55B",X"84B26A",X"4E6B35",X"000B05",X"B3C1C1",X"F6FBFF",X"FFFDFF",X"FFFCFF",X"FFFDFF",X"FDFEF8",X"FAFEF0",X"FFFFFF",X"FFFFFD",X"FEFEFC",X"FFFFFF",X"FDFDFF",X"FDFBFC",X"FFFEF7",X"F8F4E8",X"EA8631",X"E07B23",X"E97F27",X"E77D27",X"E57B2D",X"EB853B",X"E5853B",X"E08336",X"C57B4E",X"AE6D45",X"380B00",X"F1DBDD",X"FFFDFF",X"FFFFFA",X"FEFFF8",X"FBFCFF",X"FFF9FF",X"F1FDF1",X"F4FFFF",X"FEFCFF",X"F4F3F1",X"A6C083",X"80AA56",X"8BAF71",X"424F3D",X"010000",X"1B0000",X"A24C0F",X"F87712",X"FF760B",X"FF7C12",X"E47003",X"E2975D",X"FEF8EC",X"F4FFFF",X"FDFFFA",X"FCFFFF",X"FEFDF8",X"FBFFFF",X"B1D6FF",X"0E4BBE",X"196CE2",X"0068CD",X"036FD1",X"0F67E3",X"1258DA",X"1D66CC",X"2374C3",X"203C64",X"131629",X"060000",X"B9B7BC",X"FFFDFF",X"FFFCFA",X"FFFDF8",X"FCFFFF",X"FEFFFB",X"FFFFFF",X"FFFDFE",X"FFFFFB",X"FCFDFF",X"FEFBFF",X"FFFCF4",X"F9F1CA",X"E59C33",X"F97700",X"FF831C",X"ED7A0F",X"ED7B09",X"F2923E",X"BD7447",X"4E2E21",X"150000",X"380C19",X"310000",X"E9DDE9",X"FCFFFF",X"F6FCF8",X"FFFEFF",X"FFF9FF",X"FFFDFE",X"FCFEFB",X"FAF9FE",X"FDFBFE",X"ECFCFB",X"59839C",X"245892",X"3565A5",X"3A4F7C",X"2B345F",X"060022",X"1C001F",X"3D0029",X"680040",X"8C0250",X"9D0657",X"BA0D5F",X"CD126D",X"D10B6D",X"C9056B",X"C70870",X"C2036D",X"C8006F",X"DC027A",X"D10781",X"CE017A",X"D00074",X"D0006E",X"CA0068",X"C70568",X"C5106D",X"C41570",X"AC1F63",X"90275F",X"6C2955",X"4E153E",X"461034",X"1D0118",X"000909",X"00311E",X"0B8173",X"11A48A",X"01A185",X"05A58B",X"14C2A7",X"0FC0A3",X"32B19E",X"0C4743",X"03000D",X"142320",X"78A183",X"5A9B61",X"529A50",X"55954B",X"72A266",X"597A4D",X"000800",X"080500",X"976E52",X"E28C41",X"EE7910",X"FB7B1A",X"FC7E29",X"EE721A",X"FB812B",X"9C5326",X"533334",X"260F09",X"9A863F",X"C0B22F",X"C4AC18",X"D1A619",X"D1BD20",X"CBB60B",X"D2BB31",X"513D08",X"070000",X"442F1A",X"CA803F",X"FF8328",X"FF7E20",X"EE6B10",X"F27C25",X"FC8B3D",X"F07A32",X"E86F20",X"F58323",X"E4780B",X"FD7B2F",X"F67726",X"F98D35",X"D48A3F",X"724D32",X"0B0001",X"474924",X"9BA542",X"97A313",X"A8AD1B",X"9FA20D",X"ADAD19",X"B0B221",X"D9D84A",X"C7BE33",X"D0BF33",X"B69E22",X"C5AE3C",X"A69418",X"ACA125",X"BEB13F",X"BBB12E",X"B7B638",X"979A4B",X"000105",X"D3CCD3"),
(X"FFF9FF",X"929093",X"290000",X"BC2149",X"D8012B",X"D40323",X"C90628",X"D40636",X"CF022D",X"D4032D",X"D7022E",X"D1022C",X"CC052C",X"CD062F",X"D4022F",X"DB0031",X"D50C36",X"C50029",X"BB1136",X"9C283F",X"601823",X"471218",X"492024",X"381A1A",X"190909",X"000B04",X"000C0B",X"06050A",X"424333",X"7FB57B",X"78C776",X"6EAD5C",X"72B17A",X"81B58F",X"5A796A",X"040000",X"220000",X"A45B16",X"F29722",X"F18F00",X"FF9400",X"FD8F04",X"F08909",X"F18910",X"F58B1D",X"FBA04D",X"C88D61",X"290900",X"0D0600",X"0B1431",X"00175C",X"115AB6",X"197DDB",X"0C7EE1",X"0A7DF0",X"0071F5",X"0083DB",X"0079DB",X"0277E0",X"1B75D5",X"2F6AB0",X"27456B",X"15232C",X"000501",X"050300",X"292410",X"070000",X"472138",X"9F2D73",X"D50F7E",X"E40070",X"E4036D",X"F8098A",X"DC1081",X"D80E7E",X"E3057E",X"E80181",X"E60180",X"D1107D",X"AF257B",X"40121D",X"16050D",X"071515",X"000C00",X"070200",X"2B0400",X"A06006",X"CC8312",X"FDA160",X"B37F5A",X"010206",X"164781",X"3280ED",X"2C7EE4",X"3365A4",X"18204E",X"110700",X"4C1800",X"B66200",X"FFBC92",X"FFFDDB",X"EBFFFF",X"EFFCFF",X"FFFCEC",X"FDF7FF",X"FCFFFA",X"FEFDF9",X"FFFAF9",X"FBFDF0",X"B4D5C4",X"72A07C",X"85AE62",X"7AB84D",X"7DB353",X"7EB059",X"7BB65C",X"6AAD4E",X"6BAC52",X"95C37B",X"7D9A64",X"758882",X"F1FFFF",X"FAFFFF",X"FFFDFF",X"FDF7FF",X"FFFAFE",X"FFFFFA",X"FEFFF4",X"FFFFFF",X"FFFFFD",X"FEFEFC",X"FFFFFF",X"FDFDFF",X"FDFBFC",X"FFFEF7",X"F8F4E8",X"F08C37",X"DB761E",X"E1771F",X"DE741E",X"D2681A",X"C45E14",X"AA4A00",X"9F4200",X"883E11",X"450400",X"220000",X"F9E3E5",X"FCF7FB",X"FFFFFA",X"FEFFF8",X"FAFBFF",X"FFF7FF",X"F8FFF8",X"F1FFFC",X"F7F5FF",X"FFFFFD",X"A1BB7E",X"7BA551",X"769A5C",X"000600",X"0A0907",X"290500",X"C56F32",X"FF801B",X"FE6D02",X"FF841A",X"E47003",X"DB9056",X"FDF7EB",X"F4FFFF",X"FDFFFA",X"FCFFFF",X"FEFDF8",X"F9FFFF",X"84A9DD",X"0946B9",X"1D70E6",X"016DD2",X"0064C6",X"065EDA",X"1C62E4",X"1760C6",X"0354A3",X"000F37",X"0F1225",X"090003",X"C5C3C8",X"FFFEFF",X"FFF6F4",X"FFF7F2",X"FCFFFF",X"FEFFFB",X"FFFFFF",X"FFFDFE",X"FFFFFB",X"FCFDFF",X"FFFCFF",X"FFFCF4",X"FAF2CB",X"DE952C",X"FF820A",X"FD7E17",X"FA871C",X"F48210",X"D97925",X"6E2500",X"180000",X"210208",X"4B1F2C",X"5A150E",X"EFE3EF",X"F9FDFC",X"FBFFFD",X"F6F4F5",X"FFFBFF",X"FFFCFD",X"FCFEFB",X"FDFCFF",X"FEFCFF",X"ECFCFB",X"49738C",X"00326C",X"114181",X"000633",X"000934",X"0E022A",X"3D0F40",X"762462",X"8E1B66",X"B22876",X"B51E6F",X"BF1264",X"CE136E",X"CB0567",X"C40066",X"CB0C74",X"C80973",X"C8006F",X"DA0078",X"D00680",X"CE017A",X"D00074",X"D40472",X"D40972",X"CC0A6D",X"BE0966",X"B80964",X"A6195D",X"760D45",X"380021",X"250015",X"330021",X"150010",X"284646",X"408F7C",X"249A8C",X"14A78D",X"13B397",X"12B298",X"07B59A",X"0CBDA0",X"2FAE9B",X"346F6B",X"01000B",X"4D5C59",X"5E8769",X"69AA70",X"51994F",X"5C9C52",X"6F9F63",X"80A174",X"354A37",X"040100",X"4E2509",X"DC863B",X"F37E15",X"F0700F",X"FF832E",X"FF842C",X"F07620",X"CC8356",X"523233",X"140000",X"5C4801",X"B6A825",X"CAB21E",X"D6AB1E",X"CDB91C",X"C9B409",X"D4BD33",X"8A7641",X"0C0201",X"130000",X"B66C2B",X"FB7B20",X"FF7113",X"FA771C",X"E8721B",X"EF7E30",X"FF8B43",X"F98031",X"E97717",X"EC8013",X"FF863A",X"F57625",X"E1751D",X"C67C31",X"613C21",X"090000",X"545631",X"B6C05D",X"BFCB3B",X"C4C937",X"D7DA45",X"CFCF3B",X"DADC4B",X"C4C335",X"CDC439",X"DECD41",X"DCC448",X"E9D260",X"E0CE52",X"C9BE42",X"D3C654",X"DCD24F",X"DCDB5D",X"96994A",X"040509",X"DCD5DC"),
(X"FFFCF4",X"8E9295",X"0A0000",X"7C2337",X"BE1323",X"D20019",X"D7052A",X"CF0634",X"D9022E",X"DA012C",X"DB002B",X"D90028",X"D50026",X"D50026",X"D70029",X"D9002B",X"C90126",X"D8052E",X"CE0027",X"BA001F",X"C20D2E",X"CE1235",X"C60C31",X"C11334",X"740727",X"20020A",X"0A2111",X"000700",X"67713F",X"96C67A",X"6AB45B",X"78BC67",X"62AE54",X"79BB64",X"85B977",X"578264",X"00100E",X"000100",X"87643E",X"E7AB63",X"DD8311",X"F8931F",X"FF8D12",X"FF8B05",X"FF9508",X"F28D09",X"F6A031",X"DA8D31",X"562B00",X"1D0000",X"130000",X"000004",X"14324C",X"3872A4",X"2273C2",X"1672D5",X"0074E4",X"0370E9",X"1275F7",X"0C71F7",X"0E78F2",X"1879E0",X"1560B1",X"002869",X"000935",X"000225",X"06071C",X"351628",X"8A3459",X"C12E75",X"CC1378",X"D10F82",X"E20086",X"F3028D",X"E70487",X"DE007C",X"DE0175",X"D4267F",X"942C5D",X"5B122D",X"100106",X"000702",X"002D1E",X"185A4E",X"0D3735",X"00020B",X"04000B",X"120715",X"66543C",X"433029",X"0A0007",X"2A3048",X"446181",X"3B607A",X"1F3946",X"1C222E",X"1B2036",X"100600",X"70505B",X"FBE1C8",X"FFFAFF",X"FEFEFE",X"FCFDF8",X"FFFAFF",X"FFFAFF",X"FCFFF4",X"F8FAF7",X"FFF4FF",X"FFF6F6",X"95958B",X"000800",X"8B9C89",X"97B56B",X"7AA354",X"84BC65",X"74B35A",X"79B55D",X"7BB25F",X"7AAE63",X"79AD65",X"B3C3B8",X"F5FFF7",X"F9F8F6",X"FFFCFD",X"FFFAFC",X"FFFDFD",X"FEFFFD",X"F9FFFB",X"FFFFFF",X"FFFFFD",X"FEFEFC",X"FFFFFF",X"FEFCFF",X"FDFBFC",X"FFFEF9",X"F7F5E9",X"766553",X"463521",X"2F1E0C",X"1C0B01",X"0C0000",X"070000",X"010000",X"010200",X"010500",X"4F6A3D",X"6C8C67",X"E0EBE3",X"FFFEFF",X"FCFDF5",X"FDFFF3",X"FFFFFA",X"FFF9FD",X"F7FFF3",X"F5FFFA",X"FBF8FF",X"FDFCF8",X"BBD1AA",X"708866",X"0A0E0D",X"05060A",X"1F0000",X"A54B0F",X"FF8C25",X"F87100",X"F66F04",X"F4750E",X"F27A0C",X"E48C4C",X"FFF2DD",X"F8FFFB",X"FFFCF1",X"FFFBF7",X"FFFBF8",X"DAF6FF",X"327ACF",X"006EE2",X"0371E2",X"0E70DB",X"0A64D2",X"1663D5",X"3067C1",X"1A3455",X"000400",X"151D1F",X"050100",X"76736E",X"F0FEFF",X"F3FCFF",X"FFFCFD",X"FFF8F5",X"FFFEFF",X"FEFFF8",X"FFFFFF",X"FFFDFF",X"FFFFFF",X"FCFDFF",X"FFFCFF",X"FFFDF3",X"FAF2CD",X"E19944",X"EE8200",X"EC880C",X"EA8B37",X"C17C55",X"3A2222",X"140000",X"2E0003",X"5E030A",X"940A1A",X"A00000",X"FFDBDA",X"F9FFF4",X"F3F9F7",X"FFFDFF",X"FFFEFF",X"FFFCFF",X"FAFEFF",X"FFFFFF",X"FFFCFD",X"FDFAF3",X"576160",X"000513",X"1B1227",X"35002C",X"600646",X"90145C",X"B51368",X"D31474",X"D1026C",X"D90470",X"D10068",X"DA0080",X"D60680",X"CD0778",X"CF0372",X"DC0376",X"D80072",X"C8006D",X"BD096D",X"C5016F",X"C80B71",X"C3176D",X"B8256B",X"A02D64",X"6E204A",X"3D0B2E",X"260524",X"000312",X"000D15",X"002324",X"003630",X"046458",X"0A7E6B",X"22AB91",X"0AA384",X"00A78B",X"01A487",X"1BB39A",X"1DB29C",X"0BA990",X"1AAE96",X"399789",X"456768",X"0D1216",X"000A01",X"5F8B6A",X"5C9C60",X"60AA5B",X"58A24D",X"5B9B4F",X"639C58",X"5F784E",X"040A06",X"0D0000",X"B17A53",X"FFA256",X"FF8733",X"FF8225",X"F58311",X"EB7A1E",X"F79532",X"B17342",X"1C0A0A",X"060800",X"968639",X"C1A225",X"F0D02F",X"D3A81D",X"E2B622",X"ECBE2B",X"BC9B2A",X"171300",X"000104",X"7E5748",X"E18147",X"E77709",X"FA851B",X"F27A19",X"F07F23",X"F38A2F",X"FC9133",X"F07B14",X"FC7C0F",X"E6791E",X"F37F28",X"F68A2F",X"F3A654",X"693E1E",X"110000",X"5F4B26",X"D5C150",X"D6CB17",X"D9C911",X"DDCA0B",X"DACC09",X"DCD814",X"D0CD0C",X"D5CA0E",X"D9C409",X"DACA13",X"D9C70D",X"DED000",X"CEBE00",X"D0B100",X"E9C81B",X"EBDA46",X"7A7523",X"030000",X"ECCED8"),
(X"FFFCF4",X"8F9396",X"0A0000",X"6B1226",X"C01525",X"CF0016",X"DB092E",X"CD0432",X"DC0531",X"D70029",X"D70027",X"D90028",X"D80029",X"D70028",X"D70029",X"DA012C",X"CE062B",X"D10027",X"D2042B",X"C5092A",X"BF0A2B",X"C60A2D",X"C2082D",X"C01233",X"8C1F3F",X"2F1119",X"000A00",X"59664A",X"B0BA88",X"89B96D",X"67B158",X"72B661",X"73BF65",X"70B25B",X"79AD6B",X"89B496",X"466361",X"030400",X"250200",X"AF732B",X"F39927",X"F08B17",X"FC860B",X"FF8C06",X"FF8D00",X"F48F0B",X"EC9627",X"F1A448",X"B38853",X"97744E",X"675241",X"000004",X"00142E",X"002052",X"1263B2",X"1C78DB",X"0A82F2",X"026FE8",X"0C6FF1",X"0C71F7",X"0872EC",X"1374DB",X"2671C2",X"386FB0",X"335884",X"2B3F62",X"000013",X"1B000E",X"490018",X"8C0040",X"C60D72",X"D71588",X"EE0592",X"EA0084",X"E60386",X"EA0B88",X"E4077B",X"BC0E67",X"6E0637",X"300002",X"1A0B10",X"000803",X"3D7A6B",X"62A498",X"5C8684",X"202932",X"120A19",X"060009",X"120000",X"0E0000",X"10050D",X"01071F",X"000525",X"000B25",X"000613",X"00030F",X"0E1329",X"080000",X"553540",X"FFF0D7",X"FFF5FC",X"FEFEFE",X"FEFFFA",X"FFF7FF",X"FFFCFF",X"FCFFF4",X"F9FBF8",X"FFF9FF",X"F5E5E5",X"101006",X"000700",X"1D2E1B",X"82A056",X"89B263",X"7CB45D",X"79B85F",X"7FBB63",X"7CB360",X"699D52",X"78AC64",X"D3E3D8",X"F4FEF6",X"FFFFFD",X"FFFCFD",X"FFF7F9",X"FFFDFD",X"FEFFFD",X"F8FFFA",X"FFFFFF",X"FFFFFD",X"FEFEFC",X"FFFFFF",X"FEFCFF",X"FDFBFC",X"FFFEF9",X"F7F5E9",X"1F0E00",X"0E0000",X"0F0000",X"0F0000",X"231512",X"483F40",X"4C4B49",X"4D4E49",X"8D9170",X"94AF82",X"84A47F",X"E7F2EA",X"FFFEFF",X"FCFDF5",X"FEFFF4",X"FFFDF8",X"FFFBFF",X"F4FFF0",X"F2FFF7",X"FFFDFF",X"FFFEFA",X"BCD2AB",X"455D3B",X"000403",X"000004",X"795241",X"E2884C",X"EF740D",X"FD7601",X"FE770C",X"F2730C",X"E76F01",X"E78F4F",X"FFF3DE",X"F7FFFA",X"FFFCF1",X"FFFBF7",X"FEFAF7",X"D0ECFF",X"0E56AB",X"0068DC",X"0775E6",X"0062CD",X"106AD8",X"1966D8",X"003791",X"011B3C",X"11190C",X"141C1E",X"060200",X"918E89",X"ECFAFF",X"F7FFFF",X"FFFBFC",X"FFF6F3",X"FFFEFF",X"FDFFF7",X"FFFFFF",X"FEFCFF",X"FFFFFF",X"FCFDFF",X"FFFCFF",X"FFFDF3",X"FAF2CD",X"D9913C",X"FB8F09",X"F49014",X"D47521",X"5F1A00",X"110000",X"26090D",X"400F15",X"81262D",X"B22838",X"9C0000",X"FFD4D3",X"FBFFF6",X"FBFFFF",X"FEF9FF",X"FEFDFF",X"FFFDFF",X"F8FCFD",X"FDFDFF",X"FFF9FA",X"FFFFF8",X"5C6665",X"000311",X"22192E",X"712D68",X"8B3171",X"A0246C",X"B21065",X"C10262",X"DA0B75",X"D6016D",X"D6016D",X"DB0081",X"CE0078",X"CA0475",X"CF0372",X"D5006F",X"D80072",X"D00875",X"C00C70",X"CE0A78",X"CE1177",X"BB0F65",X"9F0C52",X"7E0B42",X"4B0027",X"210012",X"170015",X"101322",X"2E454D",X"417475",X"418E88",X"339387",X"37AB98",X"10997F",X"0DA687",X"02A98D",X"00A083",X"0BA38A",X"15AA94",X"12B097",X"0CA088",X"167466",X"001819",X"000206",X"001209",X"598564",X"65A569",X"63AD5E",X"5DA752",X"69A95D",X"70A965",X"799268",X"252B27",X"0D0000",X"723B14",X"E48438",X"FF8430",X"F97A1D",X"EE7C0A",X"F28125",X"DD7B18",X"BC7E4D",X"554343",X"30321C",X"665609",X"D8B93C",X"C6A605",X"EBC035",X"C79B07",X"DCAE1B",X"C4A332",X"454114",X"000104",X"562F20",X"DF7F45",X"FD8D1F",X"F88319",X"F37B1A",X"F68529",X"E37A1F",X"F4892B",X"F37E17",X"FF8013",X"ED8025",X"ED7922",X"EB7F24",X"F5A856",X"986D4D",X"160003",X"614D28",X"EFDB6A",X"E2D723",X"E5D51D",X"D7C405",X"DFD10E",X"D2CE0A",X"D1CE0D",X"D6CB0F",X"DEC90E",X"D1C10A",X"E3D117",X"D3C500",X"DBCB00",X"D7B805",X"E2C114",X"D5C430",X"635E0C",X"040001",X"EACCD6"),
(X"FEFFF6",X"A6947E",X"100600",X"1E171E",X"501A28",X"B31F2F",X"D10117",X"D70625",X"DD002B",X"E0012D",X"DD022A",X"D50326",X"D00425",X"CC0323",X"D10123",X"D70329",X"D80028",X"DB0029",X"D70026",X"D90329",X"E4012C",X"E10027",X"CE0027",X"C11835",X"7B1733",X"34131C",X"000C00",X"537A5D",X"A0C091",X"8FB272",X"83AE66",X"7CAA62",X"7FB569",X"7AB065",X"6BA45D",X"74B978",X"63AD78",X"0B4423",X"000800",X"050003",X"755026",X"CB9648",X"E89C22",X"F19100",X"FD9502",X"FD930B",X"FF9814",X"F48A03",X"F68B17",X"FFA848",X"D18843",X"260000",X"160000",X"130D0D",X"000219",X"31365C",X"375BAF",X"3A78CF",X"1973D4",X"086EDA",X"0068D9",X"0B73E6",X"0274E4",X"007DE9",X"1580E8",X"1473E1",X"0141AD",X"000D5E",X"000125",X"00000B",X"210A1A",X"511D41",X"9E2362",X"CA277A",X"CC0D74",X"D2097D",X"D91F8C",X"871459",X"130007",X"091605",X"001604",X"057159",X"11B497",X"07C2A7",X"0EB9A6",X"18A594",X"2BA58C",X"1C8F6E",X"001709",X"001013",X"0C0816",X"090000",X"070A00",X"323900",X"393100",X"513E00",X"4D4E00",X"040000",X"7A7C6E",X"FCF3FF",X"FFFBFB",X"FFFAF1",X"FEF9F5",X"FCFFFF",X"FEF9FF",X"FEFFF3",X"F7FBFE",X"FFF7FF",X"FFE1D2",X"490A00",X"230000",X"150603",X"040700",X"80927A",X"91B784",X"72A55A",X"85BA60",X"7CAC56",X"7CAA61",X"78A469",X"F8F4E8",X"FFFBF0",X"FFFEF4",X"FFFEF6",X"FFFEFA",X"FFFEFC",X"FEFFFF",X"FCFFFF",X"FEFEFE",X"FFFFFD",X"FEFEFC",X"FFFEFF",X"FFFDFF",X"FEFCFF",X"FFFFFB",X"F6F6EC",X"55744B",X"3F5E32",X"789D69",X"749C67",X"6E9B62",X"7FB172",X"77AF64",X"8EC977",X"82B371",X"71BC61",X"5FA753",X"DDF8D7",X"FFFAFF",X"FEFCFF",X"FEFFFF",X"FFFDFF",X"FFFDFF",X"FAFCF7",X"FFFFF8",X"FFFBFB",X"FEFFFF",X"B2BBB6",X"0D0600",X"1A0000",X"703203",X"E0782F",X"F87912",X"F77F0E",X"ED7807",X"F87105",X"FF780A",X"F16F00",X"D88F66",X"FFFBE5",X"F9FFFF",X"FFFCFC",X"FEF4EB",X"F6FFFF",X"83B7F3",X"0060CD",X"1D77E5",X"0D67C7",X"1E6BBD",X"2F619C",X"1F344F",X"05080F",X"000005",X"0A0D16",X"24141E",X"110100",X"C2BAA3",X"F6F7EF",X"FFFDFF",X"FFFAFF",X"FBFAF5",X"F1FFF7",X"FEFFF8",X"FFFFFF",X"FFFDFF",X"FFFFFF",X"FEFFFF",X"FEFBFF",X"FFFCF6",X"FBF2D5",X"D4914A",X"F08A48",X"A26854",X"170D04",X"0B0000",X"2A0000",X"770411",X"A11836",X"B40B32",X"BD0F30",X"A80906",X"FFD5DF",X"FFFDFF",X"FBFAFF",X"FFFEFF",X"F7FFF8",X"FFFEFB",X"F3F7F8",X"FDFCFF",X"FFFAFF",X"FFF5FE",X"707271",X"040001",X"2A1325",X"6E2C69",X"A4267A",X"CA0674",X"DA0074",X"D80578",X"C2006A",X"CE0673",X"D90277",X"D90070",X"CD006B",X"CC0C6F",X"C30567",X"CA0D71",X"C01971",X"A22665",X"78214C",X"7E2553",X"631E3D",X"4E2A36",X"060000",X"000500",X"000600",X"101113",X"050007",X"254D4F",X"3F958A",X"1FAB91",X"0BB294",X"08AC93",X"0FAB96",X"0FAE98",X"08B298",X"11B99F",X"00987F",X"13977F",X"3DA695",X"539089",X"112627",X"000600",X"000E00",X"002703",X"588860",X"659B67",X"55924D",X"5EA151",X"579C49",X"63AA5C",X"58A057",X"729C5A",X"63794A",X"000400",X"0F0000",X"C08160",X"FC8B2D",X"EF7300",X"F68E1B",X"F87A13",X"FE7B20",X"EE8A35",X"7B5025",X"484148",X"635C42",X"C7B23D",X"CCAE00",X"C7B201",X"CBB20F",X"D7B611",X"E9C82B",X"6D6002",X"030000",X"150008",X"A87059",X"E48C44",X"E08036",X"F79149",X"EB8543",X"E78A4D",X"DB8047",X"E98551",X"F68B57",X"EF9A57",X"D87A47",X"D57D4D",X"DCA270",X"857158",X"020403",X"000800",X"BDC361",X"F2E237",X"DAC416",X"DBC10C",X"F1D71E",X"ECD81F",X"D2BF09",X"DEC813",X"DFC411",X"D2C912",X"D9D325",X"D1CB15",X"DED015",X"E1CA1A",X"DACB2A",X"AFAE44",X"2D3319",X"0F0100",X"ECC5C0"),
(X"FEFFF6",X"D9C7B1",X"4F4512",X"050005",X"2B0003",X"A20E1E",X"DB0B21",X"CD001B",X"DA0028",X"DB0028",X"DE032B",X"D80629",X"CF0324",X"D00727",X"DA0A2C",X"D8042A",X"DE022E",X"DB0029",X"D50024",X"D70127",X"E3002B",X"E20028",X"CD0026",X"B80F2C",X"62001A",X"160000",X"051F12",X"001100",X"456536",X"8DB070",X"91BC74",X"7EAC64",X"79AF63",X"81B76C",X"6EA760",X"6DB271",X"6AB47F",X"70A988",X"3D5347",X"080206",X"200000",X"9C6719",X"E69A20",X"ED8D00",X"FF9A07",X"FA9008",X"FA8F0B",X"FF950E",X"F58A16",X"E08222",X"DC934E",X"C29367",X"5C462F",X"080202",X"000015",X"03082E",X"001A6E",X"1C5AB1",X"1C76D7",X"1177E3",X"0D75E6",X"0068DB",X"0C7EEE",X"0075E1",X"0671D9",X"1B7AE8",X"2C6CD8",X"2C4D9E",X"1F2F53",X"0B0F1A",X"0E0007",X"210011",X"750039",X"9A004A",X"D5167D",X"D91084",X"C60C79",X"6A003C",X"1F0413",X"000600",X"1C5947",X"3CA890",X"23C6A9",X"02BDA2",X"13BEAB",X"24B1A0",X"3AB49B",X"3CAF8E",X"468678",X"153437",X"02000C",X"746B5A",X"BDC079",X"CCD36C",X"D8D06B",X"D9C668",X"CBCC7E",X"070300",X"C6C8BA",X"FEF5FF",X"FFF7F7",X"FFFCF3",X"FFFEFA",X"F6F9FF",X"FFFDFF",X"F6FAEB",X"FCFFFF",X"FFF8FF",X"E9BBAC",X"A5663D",X"421400",X"0B0000",X"10130C",X"000800",X"628855",X"8FC277",X"77AC52",X"7DAD57",X"81AF66",X"9FCB90",X"FCF8EC",X"FFFCF1",X"FFFEF4",X"FFFEF6",X"FFFDF9",X"FFFEFC",X"FEFFFF",X"FCFFFF",X"FEFEFE",X"FFFFFD",X"FEFEFC",X"FFFEFF",X"FFFDFF",X"FEFCFF",X"FFFFFB",X"F6F6EC",X"9DBC93",X"86A579",X"89AE7A",X"8EB681",X"8AB77E",X"7DAF70",X"7CB469",X"74AF5D",X"7EAF6D",X"66B156",X"579F4B",X"E1FCDB",X"FFFDFF",X"FCFAFF",X"F9FAFF",X"FFFDFF",X"FFFEFF",X"FEFFFB",X"F5F6EE",X"FFFDFD",X"F8F9FB",X"89928D",X"070000",X"432118",X"B57748",X"ED853C",X"F5760F",X"FA8211",X"F68110",X"F16A00",X"FF780A",X"F37101",X"DB9269",X"FAE8D2",X"F5FEFD",X"FFFDFD",X"FFFDF4",X"F3FDFF",X"6DA1DD",X"005AC7",X"247EEC",X"0963C3",X"1A67B9",X"0D3F7A",X"00031E",X"0A0D14",X"141319",X"00020B",X"0A0004",X"504033",X"F4ECD5",X"FFFFF8",X"F9F6FF",X"FFF3FC",X"FFFFFA",X"F2FFF8",X"FDFFF7",X"FFFFFF",X"FEFCFF",X"FFFFFF",X"FDFEFF",X"FDFAFF",X"FFFCF6",X"FBF2D5",X"EAA760",X"CE6826",X"3D0300",X"080000",X"1E1101",X"3E0806",X"921F2C",X"9E1533",X"B1082F",X"BB0D2E",X"A30401",X"FFD5DF",X"FFFEFF",X"FDFCFF",X"FFFEFF",X"F9FFFA",X"FDF9F6",X"FCFFFF",X"FFFEFF",X"FAEEF8",X"FFF7FF",X"A0A2A1",X"060203",X"1E0719",X"3A0035",X"95176B",X"D30F7D",X"DA0074",X"D60376",X"C90571",X"D30B78",X"DA0378",X"E6097D",X"CE006C",X"B9005C",X"CC0E70",X"C3066A",X"B9126A",X"7A003D",X"4F0023",X"4A001F",X"390013",X"180000",X"2B241E",X"535E50",X"5D695F",X"1A1B1D",X"030005",X"0C3436",X"378D82",X"1EAA90",X"00A486",X"06AA91",X"1DB9A4",X"0FAE98",X"00AA90",X"05AD93",X"16AE95",X"1B9F87",X"07705F",X"00140D",X"000F10",X"000600",X"20462F",X"669470",X"75A57D",X"588E5A",X"609D58",X"589B4B",X"509542",X"5AA153",X"569E55",X"709A58",X"73895A",X"000300",X"0B0000",X"8B4C2B",X"F48325",X"F47800",X"FB9320",X"FD7F18",X"FF8025",X"EC8833",X"A0754A",X"040004",X"544D33",X"C1AC37",X"D6B80A",X"C4AF00",X"DBC21F",X"D0AF0A",X"D9B81B",X"A5983A",X"17140B",X"351E28",X"7F4730",X"D67E36",X"DE7E34",X"EF8941",X"F48E4C",X"D27538",X"CE733A",X"E37F4B",X"D06531",X"CA7532",X"E88A57",X"CA7242",X"D49A68",X"5B472E",X"000100",X"000700",X"B6BC5A",X"EBDB30",X"DEC81A",X"E7CD18",X"E5CB12",X"F9E52C",X"F1DE28",X"EFD924",X"EBD01D",X"E4DB24",X"D1CB1D",X"D2CC16",X"D2C409",X"F5DE2E",X"D8C928",X"A6A53B",X"000500",X"4C3E31",X"FFE0DB"),
(X"FEF9FF",X"F5DE90",X"B59A0D",X"1E0D00",X"050400",X"220800",X"862829",X"B91B4E",X"BE0F2E",X"C90126",X"E0002A",X"E4002A",X"D30023",X"CD0424",X"D30627",X"D60021",X"CF082F",X"CC0429",X"CC0526",X"D50328",X"E3002B",X"E1002F",X"BB0B31",X"8D162C",X"0C0100",X"00080D",X"000619",X"000219",X"00050E",X"182917",X"6F8B62",X"8FB27C",X"82A759",X"80B366",X"7EBE70",X"6AB361",X"71B663",X"7CB86E",X"82B57C",X"3A693D",X"000400",X"050800",X"76633B",X"CD9856",X"F29E3E",X"EC830E",X"FD8D0D",X"FF9A14",X"FD9001",X"FF9414",X"FF8B1A",X"FD9122",X"EA9226",X"BA7821",X"4C2000",X"1C0000",X"1A191F",X"000209",X"223D4E",X"33678F",X"2D7AC0",X"1977D7",X"0A6FDB",X"0C70E0",X"1F6CEC",X"0B70E4",X"0473DF",X"1476E3",X"1D74DD",X"0E5AB8",X"00277C",X"00004C",X"000117",X"0D1023",X"39162E",X"692D49",X"370D25",X"0B000E",X"000B07",X"00452E",X"31B4AC",X"1EB9A9",X"05B9A0",X"00BB9C",X"03C19F",X"00BD97",X"04C79B",X"00BD8C",X"36BBA6",X"1B645D",X"000302",X"91864E",X"F7F45B",X"ECEA23",X"ECE326",X"E4D927",X"F5EC25",X"B3AD19",X"D5C9BB",X"FFFEFB",X"FFFFFD",X"FAFCF7",X"F8FEFE",X"F8FFF3",X"FFFCFF",X"FEFFFA",X"EEEFF3",X"FFF8F4",X"F0A669",X"E16F0F",X"D67227",X"7A4010",X"130000",X"180300",X"120705",X"929F81",X"87B06C",X"7EB25D",X"749C53",X"CAE1AB",X"FCFCFE",X"FDFEFF",X"FBFFFF",X"F9FFFF",X"F8FFFE",X"FCFFFF",X"FFFEFF",X"FFFCFF",X"FDFFFE",X"FFFFFD",X"FEFEFC",X"FFFEFF",X"FFFDFF",X"FDFDFF",X"FFFFFB",X"F4F7EE",X"92B772",X"82AB5F",X"80AD5A",X"81B35C",X"81B65E",X"72A94E",X"8BC561",X"74AE47",X"759E58",X"71AF4E",X"6CA348",X"E8F7D0",X"FFF9FF",X"FFFCFF",X"FCFFFF",X"FFFFFD",X"FAFDFF",X"FFF9FF",X"FFFCFA",X"F6F2F3",X"FBF8FF",X"957F81",X"2A0000",X"B86D1C",X"F27911",X"FF7100",X"FF7400",X"EB6F00",X"FC7D08",X"FF7607",X"FB791B",X"D97D32",X"A07B73",X"F9F8F3",X"F5FFFF",X"F9F9FF",X"FEFCFF",X"D3E6F5",X"598DC6",X"1965B9",X"34609F",X"253F5A",X"19182A",X"0F0015",X"0F0004",X"1A0000",X"230000",X"632900",X"A05C1F",X"D0A57A",X"FFFAE3",X"FFF9F3",X"FFF9FB",X"FFFBFF",X"FCFFFF",X"F5FFFF",X"FEFFFA",X"FFFEFF",X"FEFBFF",X"FEFEFC",X"FBFDFA",X"FDFAFF",X"FFFAFB",X"FCF0E0",X"B5848A",X"411500",X"100100",X"30000A",X"7C001B",X"B10F38",X"BE0223",X"C40225",X"BD0426",X"C90D30",X"A30207",X"FCDAE8",X"F8FFFF",X"FDFAFF",X"FFFBFC",X"F7FFF6",X"FFFCFF",X"FEFFFF",X"F6F8F7",X"FFFEFF",X"F4FDFA",X"85A782",X"527944",X"001100",X"1D1D13",X"4E122B",X"A51E63",X"D0167B",X"CD0275",X"C30070",X"D0067E",X"CC007C",X"C10866",X"BF1367",X"B7256C",X"8E225E",X"520D3C",X"280820",X"070200",X"000700",X"091200",X"2C4527",X"518054",X"5A9964",X"68A973",X"79AE80",X"446747",X"000A00",X"040007",X"295A56",X"269D89",X"02A68B",X"1AC4AA",X"13B09B",X"10A28F",X"129F8C",X"2EAC96",X"4B8881",X"2B3537",X"000903",X"000D02",X"000600",X"3E5634",X"5D935F",X"5DA961",X"569C56",X"5E9D57",X"59924B",X"6CA257",X"73AB64",X"609B5B",X"639E66",X"659E5A",X"678257",X"414743",X"2C2630",X"390600",X"DA6A28",X"FF8324",X"EC8123",X"FF8615",X"F57619",X"FF8A32",X"E87E32",X"3E0500",X"362E2C",X"858756",X"CBBD42",X"CBBA15",X"DBC91F",X"E2C915",X"C3A800",X"DDC73D",X"534600",X"0B0000",X"3D2837",X"594336",X"4D3626",X"482B1B",X"633831",X"3C050B",X"6F3649",X"451A2E",X"160009",X"190000",X"865C66",X"613246",X"6F4B57",X"342333",X"0B051F",X"040005",X"8C8269",X"AAA970",X"AAA969",X"C0B975",X"B3A461",X"BFA769",X"B29A5C",X"BCAA68",X"B6AE65",X"BBAA52",X"C3BD67",X"C6BD58",X"DAC22C",X"DAC605",X"D4D027",X"9F994D",X"0E0000",X"724929",X"FFD3B5"),
(X"FFFDFF",X"E8D183",X"E1C639",X"938257",X"070601",X"311706",X"570000",X"A20437",X"C11231",X"CF072C",X"DF0029",X"E30029",X"D80528",X"D00727",X"D40728",X"E1062C",X"CB042B",X"CF072C",X"D30C2D",X"D60429",X"E10029",X"E40232",X"BB0B31",X"7E071D",X"080000",X"0B1419",X"697E91",X"58677E",X"00030C",X"000800",X"001100",X"5A7D47",X"93B86A",X"83B669",X"64A456",X"71BA68",X"71B663",X"6CA85E",X"80B37A",X"85B488",X"535F5B",X"070A00",X"120000",X"794402",X"E08C2C",X"F48B16",X"F68606",X"F78B05",X"FF9304",X"F98808",X"F98514",X"FE9223",X"F0982C",X"E19F48",X"B98D5E",X"512F23",X"000005",X"0C151C",X"000B1C",X"00153D",X"08559B",X"1B79D9",X"0A6FDB",X"177BEB",X"0B58D8",X"0F74E8",X"0F7EEA",X"0C6EDB",X"166DD6",X"2E7AD8",X"3562B7",X"2B3283",X"09142A",X"070A1D",X"16000B",X"270007",X"2A0018",X"07000A",X"0A2D29",X"489D86",X"2BAEA6",X"0CA797",X"03B79E",X"04C5A6",X"01BF9D",X"00B38D",X"02C599",X"00C392",X"2CB19C",X"2F7871",X"000403",X"675C24",X"E6E34A",X"EDEB24",X"D7CE11",X"DBD01E",X"EEE51E",X"E1DB47",X"FCF0E2",X"FFFEFB",X"F5F5F3",X"FEFFFB",X"FBFFFF",X"F6FFF1",X"FFFDFF",X"FDFFF9",X"FEFFFF",X"FFF3EF",X"E69C5F",X"DF6D0D",X"EA863B",X"C48A5A",X"402D1F",X"0F0000",X"0D0200",X"354224",X"7BA460",X"88BC67",X"8BB36A",X"D1E8B2",X"FEFEFF",X"FEFFFF",X"FBFFFF",X"F8FFFE",X"F9FFFF",X"FCFFFF",X"FFFEFF",X"FFFCFF",X"FDFFFE",X"FFFFFD",X"FEFEFC",X"FFFEFF",X"FFFDFF",X"FDFDFF",X"FFFFFB",X"F4F7EE",X"81A661",X"93BC70",X"82AF5C",X"76A851",X"6FA44C",X"77AE53",X"649E3A",X"77B14A",X"739C56",X"74B251",X"6DA449",X"E4F3CC",X"FFF5FB",X"FFFDFF",X"FCFFFF",X"FEFEFC",X"F7FAFF",X"FFFCFF",X"FCF2F0",X"FFFEFF",X"FBF8FF",X"7C6668",X"8D5830",X"CF8433",X"F87F17",X"FC6B00",X"FF7800",X"FB7F05",X"FB7C07",X"FF7607",X"FF7D1F",X"BD6116",X"926D65",X"FAF9F4",X"F2FFFF",X"FCFCFF",X"FFFEFF",X"C7DAE9",X"134780",X"0D59AD",X"0B3776",X"001631",X"000011",X"0C0012",X"19050E",X"6D5346",X"A0744F",X"BF8546",X"D18D50",X"F9CEA3",X"FFF6DF",X"FFFAF4",X"FFFDFF",X"FFFBFF",X"F9FDFF",X"F6FFFF",X"FEFFFA",X"FFFEFF",X"FEFBFF",X"FEFEFC",X"FBFDFA",X"FDFAFF",X"FFFBFC",X"FDF1E1",X"6D3C42",X"220000",X"281912",X"4D1727",X"951634",X"B00E37",X"C10526",X"BF0020",X"BB0224",X"CD1134",X"A30207",X"FCDAE8",X"F8FFFF",X"FDFAFF",X"FFFBFC",X"F6FFF5",X"FFFCFF",X"F9FAFE",X"FBFDFC",X"FFFEFF",X"F9FFFF",X"88AA85",X"789F6A",X"3C5434",X"020200",X"490D26",X"8A0348",X"BE0469",X"D90E81",X"CE077B",X"CA0078",X"D20482",X"CE1573",X"BE1266",X"930148",X"640034",X"3A0024",X"14000C",X"433E3A",X"636D54",X"79826F",X"6F886A",X"92C195",X"71B07B",X"54955F",X"609567",X"769979",X"314732",X"040007",X"001814",X"118874",X"0FB398",X"02AC92",X"0EAB96",X"21B3A0",X"19A693",X"05836D",X"002C25",X"030D0F",X"000600",X"000600",X"5C6854",X"819977",X"689E6A",X"4B974F",X"63A963",X"51904A",X"5B944D",X"7DB368",X"74AC65",X"538E4E",X"71AC74",X"6BA460",X"5B764B",X"222824",X"2D2731",X"824F3C",X"EC7C3A",X"FF892A",X"F68B2D",X"F97A09",X"ED6E11",X"F77B23",X"EB8135",X"8A5134",X"100806",X"303201",X"B0A227",X"BFAE09",X"C3B107",X"D8BF0B",X"CCB100",X"D0BA30",X"B1A45E",X"0C0000",X"382332",X"150000",X"120000",X"190000",X"1F0000",X"5D262C",X"3F0619",X"390E22",X"260719",X"55392B",X"250005",X"300115",X"180000",X"231222",X"07011B",X"3F3840",X"0E0400",X"0C0B00",X"0A0900",X"2C2500",X"433400",X"3C2400",X"180000",X"210F00",X"1F1700",X"312000",X"3E3800",X"635A00",X"CFB721",X"DBC706",X"DDD930",X"625C10",X"291419",X"896040",X"FACBAD"),
(X"FFF8EC",X"F1DE7F",X"EEC507",X"F7BD2E",X"927D12",X"000E00",X"100C00",X"480816",X"7C1824",X"A72237",X"C61436",X"D0012B",X"DA032C",X"D40028",X"D20024",X"DC042D",X"EA002B",X"E4012E",X"DB072D",X"D70127",X"DE002A",X"D40C3A",X"85182F",X"230F0E",X"000207",X"187374",X"38D7DB",X"3FD2E6",X"04667F",X"00101E",X"00070B",X"050004",X"335031",X"88AE7B",X"8BB96E",X"78AA53",X"7BAD58",X"7BAE61",X"74AE61",X"76B767",X"6BB081",X"547B60",X"121413",X"0D0005",X"311814",X"AF8A60",X"E1A44B",X"EA971F",X"F49110",X"ED8709",X"FE9516",X"FE960F",X"F59107",X"E78B06",X"FAA330",X"EF9936",X"BB7434",X"4C1600",X"180000",X"15060D",X"110C12",X"212E3E",X"3A5F8C",X"366BB7",X"2683C8",X"1475C4",X"0D70CE",X"0D74DD",X"0473DF",X"0071DD",X"0074E1",X"0A7AE8",X"1F68CF",X"003483",X"001C54",X"000023",X"070E1E",X"000107",X"2D3D3A",X"5C8B7B",X"3FAFA1",X"37B8A2",X"1FB89A",X"08B391",X"0DBEA1",X"08B8A3",X"0AB4A7",X"08AFA8",X"24CCB3",X"2C8776",X"000500",X"66540A",X"EDE230",X"F4EC0D",X"D8D100",X"E5E513",X"EEDF00",X"F8DF8D",X"FFF6E3",X"FAF8FF",X"F9FFFF",X"F5FCFF",X"FBFFFA",X"F9FFF0",X"FFFEFF",X"FAFEFF",X"FFFBFD",X"FFDDB8",X"DB7812",X"FF7C04",X"EC6803",X"E87C1A",X"D06F22",X"601500",X"230000",X"190000",X"160704",X"6D6862",X"A6ADA5",X"E7FBF2",X"FAFFFF",X"FBFFFF",X"F8FFFF",X"F8FFFF",X"FBFFFF",X"FEFFFF",X"FFFEFF",X"FFFEFF",X"FDFFFE",X"FFFFFD",X"FFFEFC",X"FFFEFF",X"FFFDFF",X"FDFCFF",X"FEFFFD",X"F2F8EE",X"73B261",X"67A952",X"71B65B",X"61A74E",X"5FA753",X"6AAE61",X"65A85B",X"72B266",X"7DAA69",X"78A85C",X"719452",X"EAF3D8",X"FFFDFD",X"FFFFFB",X"FBFEF3",X"FEFFF5",X"F8FFFF",X"FFF6FB",X"FFFBFF",X"FDFEFF",X"FFF4E7",X"C78054",X"E3731F",X"FA8011",X"FA7202",X"FF7000",X"FC7100",X"FD7E09",X"E96B05",X"ED792E",X"D28559",X"381801",X"A4999D",X"FCFEFF",X"F5FFFF",X"FDFEFF",X"F6F1F8",X"B5B9B8",X"000300",X"251D28",X"110000",X"150000",X"200000",X"6C2F10",X"B96D15",X"F1921A",X"FD881F",X"FF8C2E",X"D57600",X"FBCE97",X"FFFCFF",X"FEFEFF",X"FBFBFB",X"F8FFFF",X"FAFDFF",X"FFF9FF",X"FEFFFB",X"FFFEFF",X"FEFCFF",X"FFFFFA",X"FCFFF8",X"FEFBFF",X"FFFAFF",X"FDEFEE",X"343841",X"4E0000",X"800A20",X"9C0224",X"C40725",X"C10024",X"CD022F",X"B80034",X"AD0715",X"BA192B",X"900701",X"F7DEE4",X"F7FFFE",X"FEFDFB",X"FFFDFD",X"F7FFFB",X"FFFDFF",X"F8FBFF",X"FEFFFB",X"FDFDF5",X"F1FFEE",X"8BBC7A",X"5A9A39",X"6DA358",X"0B2E06",X"1B291C",X"1D0017",X"7F245F",X"AE1A66",X"C01865",X"B61B5F",X"AE2865",X"842E5B",X"420213",X"2E0400",X"290500",X"2A0500",X"220500",X"332B1E",X"85937A",X"70AB73",X"5E9A5E",X"619F5E",X"6EAD67",X"609F59",X"67A260",X"679D61",X"4D8048",X"091706",X"111811",X"092121",X"3F8A83",X"2AAB95",X"1AA68B",X"389E89",X"285D53",X"000600",X"040700",X"000700",X"0B300E",X"5F8E62",X"6D9465",X"699B5E",X"5EA85B",X"59A050",X"5A9E53",X"8BC882",X"679B59",X"5C8A4C",X"6D945F",X"779770",X"90AD8F",X"80947B",X"070000",X"180000",X"67351A",X"D28149",X"FF8F4B",X"FF8535",X"F78B28",X"EC7B1B",X"F1983A",X"E58D46",X"EA8B53",X"AE6F43",X"0A0000",X"020400",X"82721B",X"CBA924",X"BF9A03",X"CDA801",X"CCAD04",X"C7AC07",X"D7C138",X"675A14",X"040100",X"1D131E",X"4D1D37",X"6B0B39",X"740039",X"B93684",X"CB4A9D",X"7D004C",X"990E61",X"A11369",X"970768",X"A91E83",X"B63995",X"60004B",X"400039",X"460944",X"4A1647",X"240012",X"290018",X"280017",X"24000C",X"2D000C",X"3E0020",X"250314",X"060000",X"0C0112",X"021000",X"050C00",X"A7931A",X"EEE22A",X"BEC63C",X"4A411A",X"643136",X"C17A5A",X"FFCEA8"),
(X"FFF9ED",X"EDDA7B",X"E7BE00",X"FBC132",X"D8C358",X"546926",X"120E00",X"2E0000",X"500000",X"8F0A1F",X"C10F31",X"D1022C",X"DB042D",X"D8042C",X"D20024",X"D50026",X"EA002B",X"E0002A",X"D30025",X"D40024",X"E1002D",X"D10937",X"770A21",X"120000",X"00070C",X"45A0A1",X"3AD9DD",X"29BCD0",X"5CBED7",X"3B7583",X"001418",X"070206",X"000C00",X"002000",X"76A459",X"91C36C",X"82B45F",X"7AAD60",X"6FA95C",X"78B969",X"6EB384",X"8FB69B",X"6F7170",X"0F0007",X"140000",X"220000",X"A96C13",X"EE9B23",X"F89514",X"EE880A",X"FF9617",X"F9910A",X"F8940A",X"FCA01B",X"DF8815",X"EB9532",X"E59E5E",X"BB8561",X"755351",X"0A0002",X"09040A",X"000919",X"000B38",X"002672",X"0764A9",X"1475C4",X"187BD9",X"0B72DB",X"0271DD",X"047AE6",X"0478E5",X"006DDB",X"2069D0",X"2A73C2",X"39629A",X"343E61",X"000010",X"040B11",X"000E0B",X"001B0B",X"017163",X"13947E",X"24BD9F",X"1DC8A6",X"14C5A8",X"02B29D",X"04AEA1",X"0BB2AB",X"19C1A8",X"25806F",X"000700",X"827026",X"F3E836",X"E9E102",X"ECE510",X"F3F321",X"F1E203",X"FCE391",X"FFF7E4",X"FFFDFF",X"F5FCFF",X"F9FFFF",X"F7FCF6",X"FCFFF3",X"FEFAFB",X"FCFFFF",X"F6F0F2",X"FDD1AC",X"CC6903",X"FF7700",X"FF7C17",X"E27614",X"DA792C",X"CF844D",X"83553D",X"120000",X"30211E",X"050000",X"7D847C",X"F2FFFD",X"F9FEFF",X"FAFFFF",X"F8FFFF",X"F8FFFF",X"FBFFFF",X"FEFFFF",X"FFFEFF",X"FFFEFF",X"FDFFFE",X"FFFFFD",X"FFFEFC",X"FFFEFF",X"FFFDFF",X"FDFCFF",X"FEFFFD",X"F2F8EE",X"84C372",X"66A851",X"71B65B",X"6FB55C",X"6BB35F",X"65A95C",X"72B568",X"79B96D",X"7CA968",X"7FAF63",X"7C9F5D",X"F0F9DE",X"FFFDFD",X"FEFDF9",X"FCFFF4",X"FFFFF6",X"F6FFFF",X"FFFCFF",X"FFF9FD",X"F8F9FB",X"FFF6E9",X"E19A6E",X"DD6D19",X"F97F10",X"FB7303",X"FF7301",X"FF7803",X"F87904",X"FD7F19",X"F9853A",X"A25529",X"190000",X"D1C6CA",X"FBFDFF",X"F0FBFD",X"FEFFFF",X"FFFDFF",X"606463",X"030A03",X"040007",X"1E0606",X"674D36",X"9C715E",X"CD9071",X"DE923A",X"EB8C14",X"F47F16",X"F87618",X"F3941C",X"FFDEA7",X"FFFCFF",X"FDFDFF",X"F9F9F9",X"F9FFFF",X"FCFFFF",X"FFF9FF",X"FEFFFB",X"FFFEFF",X"FEFCFF",X"FFFFFA",X"FDFFF9",X"FEFBFF",X"FFFBFF",X"FDEFEE",X"4A4E57",X"530501",X"AD374D",X"C42A4C",X"B80019",X"C9002C",X"C60028",X"BC0438",X"B50F1D",X"B71628",X"880000",X"FBE2E8",X"F8FFFF",X"FEFDFB",X"FFFDFD",X"F6FFFA",X"FFFDFF",X"F8FBFF",X"FEFFFB",X"FFFFF8",X"EDFBEA",X"78A967",X"65A544",X"6AA055",X"698C64",X"000600",X"280A22",X"560036",X"AD1965",X"C11966",X"A4094D",X"920C49",X"5D0734",X"370008",X"2E0400",X"926E58",X"A17C6C",X"150000",X"070000",X"324027",X"5D9860",X"639F63",X"559352",X"65A45E",X"62A15B",X"6DA866",X"699F63",X"70A36B",X"4C5A49",X"000300",X"001313",X"18635C",X"2AAB95",X"17A388",X"00503B",X"001107",X"000500",X"090C03",X"434F3B",X"7FA482",X"7AA97D",X"769D6E",X"6D9F62",X"58A255",X"60A757",X"66AA5F",X"73B06A",X"699D5B",X"709E60",X"7CA36E",X"6C8C65",X"335032",X"1A2E15",X"0D0206",X"58353C",X"B8866B",X"E4935B",X"F07935",X"FF8939",X"F38724",X"ED7C1C",X"E2892B",X"F8A059",X"CF7038",X"662700",X"2F2219",X"010300",X"695902",X"DAB833",X"CCA710",X"CCA700",X"CBAC03",X"D1B611",X"BEA81F",X"A49751",X"0B0801",X"080009",X"50203A",X"8D2D5B",X"9D2062",X"AE2B79",X"C03F92",X"B12B80",X"AB2073",X"A3156B",X"A41475",X"A51A7F",X"B13490",X"811C6C",X"702369",X"5D205B",X"7A4677",X"692F57",X"512040",X"50223F",X"5C2344",X"732D52",X"6E2E50",X"3A1829",X"544B4E",X"372C3D",X"000600",X"69703C",X"D3BF46",X"D8CC14",X"B5BD33",X"1D1400",X"612E33",X"C27B5B",X"FFCAA4"),
(X"FFFFEF",X"EBD774",X"E8C400",X"FED018",X"E9C515",X"E6CA38",X"937D18",X"170400",X"0D0100",X"1B0A00",X"3E1911",X"6D2123",X"991C2C",X"B41531",X"C01633",X"C41A37",X"BD112B",X"D10327",X"DD0023",X"D50328",X"BC1330",X"87162A",X"380B12",X"000300",X"0B6C72",X"25D5D2",X"02E4E3",X"08D3E2",X"16CCDA",X"24D8D9",X"1CB5B3",X"0B737E",X"000820",X"000815",X"030500",X"5D674E",X"87A87D",X"81B77B",X"76B36D",X"70AD5F",X"72B85F",X"71B15B",X"91C67E",X"487242",X"000A00",X"000700",X"130A00",X"513D24",X"C68A58",X"E6A251",X"E28C15",X"F9910A",X"FF8D09",X"FF8F0E",X"FF8E0A",X"FF990A",X"F78600",X"FF9918",X"EF972D",X"C77B2F",X"925327",X"1F0000",X"0D0000",X"0C0D05",X"00050C",X"2A2C52",X"45569C",X"2F6FC6",X"1275D2",X"086BD1",X"0D69D6",X"1872E4",X"0071EE",X"0D6BE9",X"1978EC",X"2581E8",X"0F52AD",X"00246A",X"000733",X"000326",X"010000",X"040E0D",X"264945",X"42857C",X"46AFA0",X"31B79F",X"24B99B",X"18B393",X"24C2A9",X"348974",X"000600",X"75692D",X"E6DD42",X"ECDB0F",X"F9DF10",X"E9D300",X"E9DD0B",X"FEF693",X"FEFFFF",X"F2FFF6",X"F8FFE6",X"FFFBFF",X"FFF8FF",X"FFFBFF",X"FFFEF8",X"F8FDFF",X"FFFBFB",X"FFC288",X"E57200",X"FF7304",X"FF7518",X"FF7100",X"FF7303",X"F37006",X"EE862F",X"914A14",X"2D0700",X"0F0000",X"89807B",X"FFFEF3",X"FFFCF7",X"FFFDFA",X"FFFDFD",X"FFFCFF",X"FFFDFF",X"FFFEFD",X"FFFFFD",X"FFFFFB",X"FDFFFE",X"FFFFFD",X"FFFEFC",X"FFFEFF",X"FFFDFF",X"FDFCFF",X"FEFFFD",X"F2F8EE",X"6F9D5D",X"7EB067",X"639A47",X"79B15A",X"75AC58",X"82B664",X"669545",X"93BF70",X"6CB55C",X"7EB967",X"7DA26C",X"E6F7E5",X"F7FDFB",X"FDFFFA",X"FFFFFF",X"FFFCFF",X"F8FFFA",X"FEF6F3",X"FAF8FD",X"F8FFFF",X"F9DFAC",X"F58B25",X"FF7204",X"FF660F",X"FF7C10",X"ED6907",X"F17618",X"EA7C23",X"D67D41",X"804533",X"2D1012",X"070000",X"E0DCD9",X"FFFBFF",X"F8F8EE",X"FFFCE9",X"F2DFE5",X"261000",X"754600",X"B85E22",X"CA7439",X"EB8A19",X"FF8D0F",X"FF8312",X"F37C00",X"F98C09",X"FF911B",X"F18103",X"EEA45B",X"FFEFDB",X"F2FFFF",X"FFFDFF",X"FFFCF6",X"F4F9FC",X"F8FFFF",X"FFFEF3",X"FCFEFB",X"FFFEFF",X"FEFCFF",X"FFFFF8",X"FDFFF7",X"FEFBFF",X"FFF9FF",X"FCEDF4",X"873F4B",X"850000",X"D22D4D",X"E83263",X"B6002B",X"A80429",X"B70E21",X"B50919",X"AE1534",X"6C202D",X"350A00",X"F0E6F1",X"FFF7FD",X"FFFAF6",X"F9FFFD",X"FAFBFF",X"FDFFFE",X"F8FDFF",X"FFFFFB",X"FBF0F4",X"FFFEFF",X"85A97D",X"5E9248",X"6E996E",X"80A675",X"597D63",X"000A0E",X"281630",X"4D1636",X"5D1932",X"2A0001",X"160000",X"250000",X"884211",X"D77224",X"FA8C35",X"DB833C",X"4F1F00",X"070000",X"02131B",X"6B985F",X"6DA161",X"5D9A54",X"60A457",X"63AA5A",X"5EA152",X"659F53",X"6EA35B",X"6E946B",X"102D0F",X"000900",X"051719",X"455D5F",X"253B39",X"000500",X"050800",X"0A2B0E",X"547E58",X"7AB380",X"69AD72",X"539859",X"70B16F",X"65A75D",X"5BA04D",X"669C51",X"82B975",X"62985A",X"74A76E",X"6F9967",X"56704B",X"000500",X"070700",X"190000",X"683812",X"CD804A",X"F48939",X"F47A17",X"FC801E",X"EE7725",X"E97730",X"F3823C",X"D5925B",X"A48B62",X"332717",X"070002",X"080100",X"917D24",X"DAAD36",X"C6AC0D",X"D5AD10",X"C99D08",X"E0BE27",X"D3B20B",X"DAB409",X"CAAC26",X"7B6D15",X"000911",X"110015",X"6E1A55",X"A41370",X"BE0177",X"C50071",X"CD0170",X"C80264",X"CB0A7D",X"C8077A",X"D20C83",X"C60072",X"D60E7B",X"CE1072",X"CB1C7B",X"CA2486",X"D31380",X"BA0E74",X"B11171",X"B81477",X"BD127A",X"AF1671",X"8C2366",X"8A4B78",X"351C32",X"3E4A26",X"BBBD7C",X"F1D065",X"F2DC4B",X"A4AB5B",X"0B0000",X"B8765C",X"C97B65",X"FFD5B3"),
(X"FCFFEC",X"EEDA77",X"F0CC00",X"F1C30B",X"E3BF0F",X"E3C735",X"E7D16C",X"B3A068",X"3A2E22",X"0D0000",X"1B0000",X"4E0204",X"79000C",X"950012",X"B10724",X"BE1431",X"C31731",X"D90B2F",X"E5032B",X"DD0B30",X"B9102D",X"720115",X"240000",X"000300",X"3A9BA1",X"27D7D4",X"00DBDA",X"0DD8E7",X"19CFDD",X"1CD0D1",X"32CBC9",X"4BB3BE",X"405C74",X"000512",X"020400",X"000700",X"2F5025",X"79AF73",X"73B06A",X"75B264",X"68AE55",X"75B55F",X"70A55D",X"97C191",X"6F8872",X"000500",X"080000",X"140000",X"3D0100",X"965201",X"E58F18",X"FF9912",X"FD8804",X"FF900F",X"FB8A06",X"F58C00",X"FF9205",X"FC9514",X"E99127",X"E5994D",X"E3A478",X"936A54",X"342319",X"000100",X"00050C",X"000026",X"00054B",X"003087",X"086BC8",X"1A7DE3",X"1571DE",X"126CDE",X"0173F0",X"0967E5",X"1372E6",X"106CD3",X"2E71CC",X"3469AF",X"254E7A",X"142144",X"050402",X"000302",X"000B07",X"001D14",X"006758",X"0D937B",X"11A688",X"20BB9B",X"2BC9B0",X"3F947F",X"000400",X"564A0E",X"DAD136",X"F9E81C",X"FEE415",X"F2DC00",X"EDE10F",X"FFFF9F",X"F3F4F8",X"F7FFFB",X"FCFFEA",X"FFFDFF",X"FFF1FF",X"FFFBFF",X"FFFEF8",X"F5FAFE",X"FDF1F1",X"E6A56B",X"E67300",X"FF7A0B",X"FF7114",X"FF7402",X"FE6E00",X"FF7F15",X"D87019",X"D18A54",X"825C47",X"1C0A08",X"D0C7C2",X"FFFAEF",X"FFFCF7",X"FFFDFA",X"FFFDFD",X"FFFCFF",X"FFFDFF",X"FFFEFD",X"FFFFFD",X"FEFFFA",X"FDFFFE",X"FFFFFD",X"FFFEFC",X"FFFEFF",X"FFFDFF",X"FDFCFF",X"FEFFFD",X"F2F8EE",X"87B575",X"6FA158",X"88BF6C",X"83BB64",X"7EB561",X"8ABE6C",X"84B363",X"7EAA5B",X"7DC66D",X"74AF5D",X"658A54",X"DDEEDC",X"FBFFFF",X"FEFFFB",X"FBFBFB",X"FFF9FF",X"F7FFF9",X"FFFDFA",X"FDFBFF",X"F3FEFA",X"EFD5A2",X"E17711",X"FF7204",X"FF650E",X"FA7206",X"FE7A18",X"FB8022",X"ED7F26",X"9E4509",X"2D0000",X"3A1D1F",X"060000",X"D6D2CF",X"FFFCFF",X"FAFAF0",X"FFFDEA",X"FFF2F8",X"9E8870",X"C5964E",X"EC9256",X"E58F54",X"EC8B1A",X"FC8608",X"FB7C0B",X"FD8606",X"FE910E",X"F58610",X"F18103",X"F4AA61",X"FFFCE8",X"F0FDFF",X"FBF8FF",X"FFFCF6",X"F7FCFF",X"F9FFFF",X"FFFBF0",X"FBFDFA",X"FEFDFF",X"FEFCFF",X"FFFFF8",X"FDFFF7",X"FEFBFF",X"FFF8FF",X"FCEDF4",X"904854",X"900604",X"B10C2C",X"B1002C",X"BE0733",X"A70328",X"AE0518",X"BE1222",X"A50C2B",X"550916",X"200000",X"EAE0EB",X"FFF6FC",X"FCF7F3",X"F9FFFD",X"FCFDFF",X"FCFEFD",X"FBFFFF",X"FDFCF8",X"FFF9FD",X"FAF9FE",X"92B68A",X"5F9349",X"75A075",X"789E6D",X"769A80",X"0F2226",X"22102A",X"2B0014",X"330008",X"300007",X"644845",X"A4765F",X"D08A59",X"EE893B",X"EE8029",X"DB833C",X"A3734F",X"060000",X"00040C",X"5C8950",X"7BAF6F",X"609D57",X"519548",X"5BA252",X"68AB5C",X"659F53",X"679C54",X"769C73",X"456244",X"000A00",X"000F11",X"000A0C",X"000907",X"000C03",X"35382D",X"7A9B7E",X"79A37D",X"669F6C",X"4F9358",X"5FA465",X"5FA05E",X"62A45A",X"5CA14E",X"689E53",X"619854",X"74AA6C",X"669960",X"37612F",X"000C00",X"010A00",X"010100",X"80623E",X"BE8E68",X"D58852",X"E67B2B",X"FC821F",X"FF8725",X"F57E2C",X"F6843D",X"FE8D47",X"A9662F",X"160000",X"0A0000",X"1E1319",X"817A5E",X"BDA950",X"D9AC35",X"C0A607",X"CCA407",X"D8AC17",X"D5B31C",X"C7A600",X"CAA400",X"CFB12B",X"978931",X"00030B",X"4A314E",X"76225D",X"AC1B78",X"CB0E84",X"CF027B",X"CE0271",X"D71173",X"C40376",X"C70679",X"CA047B",X"D0067C",X"C9016E",X"CD0F71",X"C81978",X"C11B7D",X"C80875",X"C0147A",X"B31373",X"BB177A",X"B2076F",X"A70E69",X"9A3174",X"370025",X"10000D",X"414D29",X"A7A968",X"A7861B",X"B29C0B",X"6F7626",X"0D0000",X"96543A",X"D1836D",X"FFD6B4"),
(X"FFF7FD",X"DDD37E",X"E9CD08",X"E8D316",X"F3CA00",X"DCC304",X"E6C200",X"F3D221",X"DABC2A",X"9D8100",X"6E5600",X"0F0200",X"0B0600",X"0D0600",X"241414",X"2F190E",X"561422",X"54192D",X"691B17",X"752B2A",X"6D212B",X"411224",X"000902",X"0B7A71",X"25DED8",X"00CBC6",X"00D6D7",X"05DEE3",X"0CD8E1",X"0CD1DA",X"05CAD3",X"0DD3DE",X"26D8E2",X"149CAC",X"00233A",X"00091C",X"000204",X"14200C",X"768B64",X"A2BD8A",X"79A766",X"7CB066",X"73B460",X"6FBB61",X"71BB6C",X"639E64",X"3C5D3E",X"000800",X"080B12",X"030106",X"1E1007",X"A07D57",X"DF9D51",X"F1942A",X"F58809",X"FF910B",X"F59711",X"F58D06",X"FF930C",X"FC8300",X"FE8D13",X"FFA337",X"DE852B",X"C97626",X"581D00",X"250000",X"100000",X"0B0B03",X"00020B",X"243C58",X"345C90",X"3668AF",X"2977C1",X"0E6BCB",X"016BE5",X"0875F6",X"0B6FE7",X"0F6EDA",X"197BE6",X"0E76E5",X"025CAA",X"003983",X"000D4E",X"000738",X"00001B",X"00000D",X"132529",X"1E3E3D",X"507E74",X"436360",X"010602",X"544A2F",X"DAC785",X"F8E177",X"E8DF54",X"F7EE53",X"EBE587",X"FFF7C4",X"FFF6F6",X"FFF9FF",X"FDFBFF",X"FDFEFF",X"FEFFFD",X"FCFDFF",X"FBFEFF",X"FFFFFB",X"FFE4ED",X"CB8B4D",X"E27000",X"F97800",X"FF7A09",X"FF7304",X"F57619",X"FF7401",X"FC7710",X"F07819",X"FF7B12",X"B7631D",X"FAEDDA",X"FFFFF1",X"FDFBFE",X"FFFCFF",X"FFFEFF",X"FFFEFF",X"FFFEFD",X"FFFDFC",X"FFFEFB",X"FFFEFB",X"FBFEFF",X"FFFFFF",X"FFFCF9",X"FFFEFA",X"FEFDFB",X"FCFEFD",X"FEFEFE",X"F3F2EE",X"99A69C",X"85995C",X"95A487",X"829575",X"728774",X"728B6E",X"738869",X"70805C",X"677262",X"393C2B",X"060100",X"ECE6D8",X"FEFFF7",X"F9FFFF",X"F7FBFC",X"FFFFFB",X"FFF1FF",X"F7FFFD",X"E8FFF0",X"FFFCE0",X"FFB770",X"E46902",X"FF7B0E",X"F47D09",X"FF7B12",X"E17A15",X"CF9354",X"795942",X"261207",X"1C0E00",X"0F0300",X"5D5540",X"F1E7E6",X"F8FFF5",X"FFF9FF",X"FCFAE3",X"FDDEA8",X"F89118",X"EF8702",X"FE8E0E",X"FF8613",X"FF8810",X"FC8505",X"FE8503",X"F87D00",X"FF8E12",X"FF9520",X"E5800C",X"E3CAA2",X"FFF4E0",X"FFFCFB",X"FBFFFF",X"FBFFFF",X"FBFDF8",X"FFFEFF",X"FFFBFF",X"FFF8FF",X"FFFCFF",X"F9FEFA",X"F8FFFC",X"FAFFFC",X"FFFFFD",X"FFFAFE",X"FCE8F1",X"9A3E53",X"B20A23",X"BD1320",X"B40017",X"C20325",X"A90D23",X"9D172F",X"7A0F2D",X"2E0817",X"1E150C",X"000500",X"ECEAED",X"FFFAFF",X"F7F6F4",X"F9FFF9",X"FCFFFF",X"FFFCF6",X"FFFCFF",X"FFFEFF",X"FBFCFF",X"F5FFFE",X"89A572",X"6B9541",X"719C64",X"819768",X"50624A",X"00030B",X"00051F",X"120D23",X"160000",X"6D3A29",X"D89376",X"FF8735",X"F87E1B",X"F47D05",X"FC8100",X"FF8308",X"E6791A",X"6E3000",X"0E0000",X"2C2218",X"86A792",X"5B9E75",X"609D61",X"6CA055",X"5C9949",X"5CA053",X"61A35C",X"5FA157",X"6B995B",X"394D2A",X"010400",X"0E121B",X"000805",X"326141",X"61A067",X"6B9F5F",X"659C58",X"639C55",X"66A35E",X"64A064",X"639D62",X"6CA362",X"619650",X"6EA65F",X"8FAF7E",X"6D7162",X"201B21",X"060108",X"120000",X"2E0000",X"B4623C",X"F99349",X"F98B2A",X"FA8013",X"FD7C14",X"F27A19",X"E4822B",X"EAA16A",X"B77D69",X"836766",X"070000",X"2D3015",X"322600",X"B68B2D",X"E2AB2C",X"E1B820",X"BEAD08",X"D5BA0B",X"C2A000",X"E4BB21",X"D3A804",X"DBB001",X"D5AF04",X"C6A615",X"CFB23A",X"80701B",X"3D3623",X"4E3150",X"771359",X"C51A82",X"C1006A",X"C60A6B",X"C21277",X"C1046B",X"C9066F",X"D20874",X"CE0470",X"C90873",X"B9006C",X"C6107F",X"D51E90",X"CB0387",X"D91291",X"D90484",X"D60076",X"B60369",X"953A77",X"2B1931",X"000407",X"060A13",X"00010A",X"01050E",X"000307",X"000409",X"000309",X"11141D",X"554D5C",X"3C3D38",X"FBD4D7"),
(X"FFF8FE",X"E4DA85",X"E9CD08",X"E3CE11",X"F3CA00",X"E4CB0C",X"EFCB00",X"EECD1C",X"E5C735",X"E3C740",X"DEC66C",X"7F723E",X"433E16",X"100900",X"0C0000",X"110000",X"330000",X"270000",X"400000",X"490000",X"440002",X"360719",X"000500",X"29988F",X"27E0DA",X"00CAC5",X"00D9DA",X"03DCE1",X"00CCD5",X"0FD4DD",X"12D7E0",X"06CCD7",X"15C7D1",X"41C9D9",X"59A4BB",X"223D50",X"000305",X"0D1905",X"000B00",X"57723F",X"82B06F",X"76AA60",X"75B662",X"6DB95F",X"6EB869",X"7CB77D",X"90B192",X"475548",X"00030A",X"010004",X"150700",X"1D0000",X"A36115",X"FB9E34",X"FF9415",X"FF8F09",X"F2940E",X"FA920B",X"FA8600",X"FF900D",X"F9880E",X"F99428",X"F69D43",X"EE9B4B",X"BB8058",X"845939",X"503E2A",X"060600",X"000710",X"000420",X"001246",X"01337A",X"07559F",X"1F7CDC",X"127CF6",X"0069EA",X"0D71E9",X"106FDB",X"0F71DC",X"0B73E2",X"247ECC",X"266EB8",X"3764A5",X"1E2E5F",X"080927",X"060815",X"000509",X"000A09",X"000F05",X"0A2A27",X"020703",X"1E1400",X"685513",X"7E6700",X"8C8300",X"BAB116",X"C5BF61",X"FFFDCA",X"FFFBFB",X"FFF5FF",X"F9F7FF",X"FEFFFF",X"FEFFFD",X"FDFEFF",X"F9FCFF",X"FFFFFB",X"FFE2EB",X"B77739",X"F38107",X"FF7E06",X"FD6A00",X"FF790A",X"EF7013",X"FF6900",X"F7720B",X"F37B1C",X"FD780F",X"D8843E",X"FFF2DF",X"FBFCEC",X"FEFCFF",X"FFFCFF",X"FFFEFF",X"FFFEFF",X"FFFEFD",X"FFFDFC",X"FFFEFB",X"FFFEFB",X"FBFEFF",X"FFFFFF",X"FFFCF9",X"FFFEFA",X"FFFEFC",X"FCFEFD",X"FEFEFE",X"F3F2EE",X"4A574D",X"324609",X"263518",X"1A2D0D",X"000900",X"001200",X"000A00",X"000C00",X"000500",X"030600",X"100B00",X"E6E0D2",X"FFFFF8",X"F6FFFE",X"FCFFFF",X"FFFFFB",X"FFF6FF",X"EEFBF4",X"EEFFF6",X"FFF5D9",X"EEA45D",X"EF740D",X"FD790C",X"EE7703",X"FF750C",X"E17A15",X"864A0B",X"220200",X"0F0000",X"50421D",X"958963",X"BAB29D",X"FFFCFB",X"FBFFF8",X"FFF7FF",X"FFFFE8",X"EBCC96",X"EC850C",X"EC8400",X"FC8C0C",X"FF901D",X"FB840C",X"FE8707",X"FF8907",X"FF8403",X"FF8B0F",X"F58813",X"E37E0A",X"F4DBB3",X"FFFCE8",X"FFFDFC",X"F8FDFF",X"FBFFFF",X"FBFDF8",X"FFFEFF",X"FFFBFF",X"FFF8FF",X"FFFCFF",X"F9FEFA",X"F8FFFC",X"FAFFFC",X"FFFFFD",X"FFF9FD",X"FBE7F0",X"A1455A",X"A70018",X"BD1320",X"C20C25",X"BC001F",X"AF1329",X"8D071F",X"5C000F",X"280211",X"080000",X"000500",X"E2E0E3",X"FFFBFF",X"FFFFFD",X"FBFFFB",X"F4F8F9",X"FFFEF8",X"FFFDFF",X"F9F7F8",X"FDFEFF",X"F3FDFC",X"8BA774",X"638D39",X"7AA56D",X"63794A",X"000800",X"000C14",X"0C132D",X"0A051B",X"170001",X"643120",X"C58063",X"FE812F",X"FA801D",X"F47D05",X"FF8504",X"FB7D02",X"F28526",X"B17342",X"0D0000",X"0C0200",X"375843",X"6EB188",X"67A468",X"609449",X"5C9949",X"67AB5E",X"62A45D",X"63A55B",X"6B995B",X"718562",X"010400",X"000009",X"425B58",X"6D9C7C",X"73B279",X"659959",X"6CA35F",X"639C55",X"68A560",X"5C985C",X"649E63",X"609756",X"689D57",X"649C55",X"50703F",X"040800",X"030004",X"060108",X"513E38",X"B17D65",X"D5835D",X"E27C32",X"F48625",X"F47A0D",X"F97810",X"F27A19",X"F29039",X"AF662F",X"410700",X"150000",X"080000",X"4B4E33",X"ACA066",X"CFA446",X"D8A122",X"D3AA12",X"C9B813",X"CDB203",X"CEAC0C",X"CCA309",X"D5AA06",X"DBB001",X"DCB60B",X"CAAA19",X"CDB038",X"B1A14C",X"231C09",X"110013",X"5F0041",X"B2076F",X"CC0675",X"EC3091",X"C11176",X"C60970",X"C5026B",X"CA006C",X"D00672",X"CF0E79",X"BA006D",X"BA0473",X"B90274",X"CE068A",X"BF0077",X"D3007E",X"E00480",X"B50268",X"892E6B",X"36243C",X"071619",X"161A23",X"0A0D16",X"000009",X"061115",X"28373C",X"0B181E",X"000009",X"332B3A",X"000100",X"EFC8CB"),
(X"FFFEDD",X"EDDA71",X"ECC200",X"ECC717",X"FAC809",X"ECC61D",X"F6CA07",X"EAC616",X"F7DB00",X"F4D40F",X"F7D51B",X"E3C819",X"E3CA3A",X"BEA62A",X"826500",X"411C00",X"0A0A00",X"2B0000",X"1D0100",X"070100",X"172434",X"060009",X"004151",X"32CBC6",X"13D8E1",X"1AD8E8",X"03C8D8",X"01DAE1",X"00E2E0",X"00D5D2",X"0BDBDD",X"0AD1D8",X"00DDE2",X"00C7CC",X"28E1E4",X"27C5C8",X"138D8E",X"00161B",X"000813",X"01000D",X"314127",X"81A17A",X"8DC087",X"71A864",X"70A55D",X"81B672",X"73B472",X"6DBC7A",X"57A358",X"325D32",X"000400",X"10060F",X"060000",X"80714A",X"BE9054",X"E39854",X"E9901C",X"E88E13",X"FFA520",X"E78E00",X"F39B06",X"FA990A",X"FD8E08",X"FF890A",X"F99E12",X"F49B25",X"EF9B43",X"9C4C11",X"430000",X"270000",X"1C0A06",X"000108",X"000109",X"314B6E",X"2F61AA",X"2769CA",X"236DD6",X"1C71DB",X"0569D8",X"0677ED",X"0469D3",X"0A73DE",X"107BE5",X"066CD1",X"0D68C5",X"0D5BAE",X"0950A0",X"002F7E",X"000D38",X"000012",X"0B0001",X"0A0004",X"17070A",X"000300",X"000600",X"060118",X"928D77",X"F6F2E9",X"FFFEFF",X"F9F9F9",X"FEFFF8",X"FFFFF3",X"FFFFFA",X"FBF9FE",X"FEFDF9",X"FFFDF5",X"DDDAED",X"381E21",X"826539",X"CE8455",X"E28537",X"E67010",X"F67E0E",X"FF7500",X"FF7805",X"FD7914",X"EC6603",X"EA9A67",X"FDF3FC",X"F8FCFF",X"FCFDFF",X"FDFEFF",X"FCFFFF",X"FCFFFF",X"FBFFFF",X"F9FFFF",X"F8FFFF",X"F8FFFF",X"FEFFFF",X"FFFEFF",X"FFFCF9",X"FFFEFB",X"FEFEFE",X"FCFEFD",X"FFFEFC",X"F7F2EE",X"2F1403",X"1C0400",X"1F0000",X"220000",X"220000",X"260000",X"400800",X"4D0E00",X"6E1E00",X"974305",X"9F5C28",X"FFE6D9",X"FFFBFF",X"FEFAFF",X"FFFEFF",X"F2FCF3",X"FCFFF6",X"F4F9F3",X"FFF9FF",X"FFDEC8",X"DE6F1E",X"F97513",X"F47D2D",X"E38638",X"936E51",X"69503C",X"080000",X"10050D",X"1C1500",X"B1AC2E",X"EDE96B",X"F4ECAD",X"FAF9FF",X"F8FFFF",X"FFF7FF",X"FFFBEB",X"E8AF82",X"F27911",X"FF7F0F",X"FF7F14",X"FC8B13",X"F5870C",X"F5870A",X"FE8D13",X"F98715",X"EF821B",X"EA8628",X"E2842A",X"FFE5D7",X"FFF9F8",X"FFFAFF",X"FBF9FF",X"FDFEFF",X"FDFDFD",X"FFFFFF",X"FCFBFF",X"F7FFFF",X"FEFFFF",X"FFFCFD",X"FFFFFF",X"FBFFFC",X"FDFFFE",X"FFF9FD",X"FDE6EE",X"C4364E",X"BE011D",X"B01123",X"9D1430",X"92213F",X"52151C",X"260704",X"0F0B08",X"000D00",X"29532D",X"6E9C77",X"DAF0E4",X"FFFEFF",X"FAFAF8",X"FBFCF7",X"FFFDFF",X"FFFFFD",X"F4F1F8",X"FFFFFF",X"F5FBF9",X"F1FFF9",X"92B386",X"75A665",X"548661",X"030102",X"000823",X"000B48",X"164B99",X"094083",X"00062B",X"040507",X"614736",X"C39154",X"EF8B2D",X"FC7605",X"F97914",X"F87D1D",X"FB7D16",X"E17E21",X"8C530E",X"0B0000",X"000205",X"6B8771",X"88AF6C",X"659D46",X"4F954D",X"64A762",X"649A46",X"669F58",X"669A5A",X"629258",X"5D8E56",X"5D9558",X"5F9D5A",X"66A763",X"52934F",X"70B878",X"51995A",X"579D5F",X"63A464",X"6FA663",X"689157",X"97B289",X"6D8064",X"243427",X"06110D",X"0D0C0A",X"140000",X"986530",X"DD8F3C",X"FB9832",X"F28619",X"E97C1F",X"ED8429",X"EF8C37",X"DE8B3F",X"C4854F",X"835A3C",X"0F0000",X"1A1309",X"4C4800",X"6C5D00",X"A68C13",X"DCC030",X"BFA506",X"C2AA02",X"CAAC00",X"DDBB04",X"CCA80A",X"DABE1F",X"D3BF20",X"BEAD07",X"CCB505",X"D1B100",X"D4AC00",X"D0A600",X"D1AA27",X"876E2E",X"080200",X"281C28",X"752B66",X"AC1670",X"B80060",X"BF006F",X"BD0678",X"C10273",X"CA0171",X"D60B77",X"D80D78",X"CB026A",X"D20971",X"CB026C",X"D4136E",X"DF2181",X"C2086D",X"B10961",X"A12B68",X"512644",X"293C4B",X"073B48",X"1E8D7C",X"1A8374",X"005E50",X"006A5A",X"2B9F8C",X"108471",X"005043",X"075E56",X"002B2A",X"C3D7DE"),
(X"FFFEDD",X"EBD86F",X"E7BD00",X"F0CB1B",X"FECC0D",X"E7C118",X"F4C805",X"EBC717",X"F0D400",X"F3D30E",X"E8C60C",X"E1C617",X"E7CE3E",X"E8D054",X"E5C860",X"CFAA66",X"A3A36D",X"CA9C5E",X"CDB18A",X"7C765E",X"182535",X"07000A",X"4A8D9D",X"38D1CC",X"05CAD3",X"24E2F2",X"0DD2E2",X"00CDD4",X"00DDDB",X"00DCD9",X"09D9DB",X"0BD2D9",X"00D9DE",X"00CDD2",X"10C9CC",X"3AD8DB",X"4BC5C6",X"3E898E",X"102C37",X"00000C",X"000800",X"012100",X"5F9259",X"81B874",X"80B56D",X"71A662",X"79BA78",X"64B371",X"6CB86D",X"86B186",X"646965",X"0C020B",X"0C0500",X"0F0000",X"6A3C00",X"9D520E",X"E78E1A",X"F79D22",X"E68B06",X"F09707",X"F09803",X"F89708",X"FE8F09",X"FF8D0E",X"EE9307",X"F69D27",X"E38F37",X"EC9C61",X"CE8864",X"7C4D3B",X"0D0000",X"01040B",X"00050D",X"000A2D",X"002069",X"1153B4",X"246ED7",X"1F74DE",X"0F73E2",X"0071E7",X"1378E2",X"0D76E1",X"046FD9",X"0F75DA",X"1B76D3",X"1866B9",X"2C73C3",X"2C6FBE",X"2A4570",X"000012",X"1A0B10",X"170711",X"150508",X"161906",X"243427",X"020014",X"BDB8A2",X"FFFFF6",X"FCFAFD",X"F9F9F9",X"FEFFF8",X"FCFEF0",X"FFFFFA",X"FFFEFF",X"FFFEFA",X"FFFCF4",X"BEBBCE",X"140000",X"190000",X"964C1D",X"DD8032",X"F68020",X"EB7303",X"FF7000",X"FE6E00",X"F97510",X"F16B08",X"FFB683",X"FFF8FF",X"F5F9FF",X"FDFEFF",X"FDFEFF",X"FCFFFF",X"FCFFFF",X"FBFFFF",X"F9FFFF",X"F7FFFF",X"F7FFFF",X"FDFEFF",X"FFFEFF",X"FFFCF9",X"FFFEFB",X"FEFEFE",X"FDFFFE",X"FFFFFD",X"F7F2EE",X"735847",X"6B5313",X"795734",X"815C32",X"8D6240",X"8D6039",X"AB7352",X"B07150",X"CA7A49",X"DA8648",X"C88551",X"FFE1D4",X"FFFBFF",X"FFFBFF",X"FFFEFF",X"F8FFF9",X"FCFFF6",X"F6FBF5",X"FFF9FF",X"FFC0AA",X"E27322",X"FE7A18",X"ED7626",X"BB5E10",X"411C00",X"170000",X"1E130F",X"070004",X"C3BC78",X"E9E466",X"E4E062",X"FFFBBC",X"FDFCFF",X"F8FFFF",X"FFFAFF",X"FFFDED",X"E7AE81",X"ED740C",X"FF8313",X"FF8217",X"F6850D",X"FD8F14",X"F28407",X"FB8A10",X"FA8816",X"EE811A",X"F28E30",X"F2943A",X"FFE8DA",X"FFF9F8",X"FFF9FF",X"FCFAFF",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FBFAFF",X"F6FFFF",X"FEFFFF",X"FFFCFD",X"FFFFFF",X"FBFFFC",X"FDFFFE",X"FFF9FD",X"FDE6EE",X"C83A52",X"BD001C",X"B11224",X"9A112D",X"7B0A28",X"340000",X"170000",X"070300",X"617663",X"87B18B",X"5F8D68",X"DEF4E8",X"FFFEFF",X"FFFFFD",X"FCFDF8",X"FDF8FE",X"FDFCFA",X"FFFDFF",X"FFFFFF",X"F9FFFD",X"F5FFFD",X"85A679",X"5B8C4B",X"043611",X"010000",X"03112C",X"1B3D7A",X"2B60AE",X"2B62A5",X"0E3055",X"050608",X"140000",X"774508",X"F38F31",X"FF7D0C",X"FF831E",X"F87D1D",X"F2740D",X"F59235",X"BA813C",X"1F100D",X"000407",X"19351F",X"8BB26F",X"6AA24B",X"5DA35B",X"589B56",X"679D49",X"5C954E",X"6CA060",X"6D9D63",X"6C9D65",X"669E61",X"70AE6B",X"66A763",X"599A56",X"559D5D",X"71B97A",X"549A5C",X"76B777",X"70A764",X"689157",X"4C673E",X"041700",X"000C00",X"000703",X"21201E",X"A88E7D",X"CC9964",X"DF913E",X"D8750F",X"FF9326",X"FF9437",X"F48B30",X"EC8934",X"C87529",X"6B2C00",X"230000",X"120000",X"171006",X"B7B36A",X"BFB053",X"C9AF36",X"BFA313",X"C0A607",X"C9B109",X"CEB000",X"D5B300",X"CDA90B",X"CDB112",X"D7C324",X"BCAB05",X"CDB606",X"DBBB08",X"DAB202",X"D7AD01",X"EAC340",X"B39A5A",X"231D0F",X"3B2F3B",X"651B56",X"A20C66",X"CB0C73",X"C60476",X"BB0476",X"C30475",X"C8006F",X"CB006C",X"CA006A",X"CA0169",X"D40B73",X"CC036D",X"C90863",X"D71979",X"BA0065",X"BA126A",X"810B48",X"2D0220",X"000615",X"3F7380",X"309F8E",X"3FA899",X"369B8D",X"2C9787",X"30A491",X"2CA08D",X"309689",X"3F968E",X"40807F",X"D5E9F0"),
(X"FCFFE4",X"EEDA79",X"EEBC03",X"F0C818",X"F4C908",X"E6BF0C",X"F5CD00",X"EDD501",X"EDCD00",X"F9CF1B",X"F4C012",X"F8C410",X"EEBF0D",X"EBC405",X"F2D00C",X"F0CB1B",X"E0E020",X"F2C208",X"F3D050",X"839160",X"000300",X"010109",X"1F4A5A",X"57B5BD",X"2BD7D9",X"14CBD3",X"12D6E4",X"06CFDF",X"00CBDA",X"05D4DE",X"00D0D7",X"08DFE4",X"06D2DD",X"03D3DD",X"07DCE4",X"00D5DB",X"0AD3DA",X"22D0DB",X"2BB8CA",X"005C75",X"000417",X"030B16",X"000200",X"3D5136",X"82AC7A",X"84BB77",X"73A95B",X"83B262",X"77A55A",X"76B268",X"79C07C",X"52965B",X"305F31",X"223B1E",X"000500",X"000100",X"422F0E",X"A8804F",X"E8A056",X"F89730",X"FA8F0F",X"FE9505",X"FF9C03",X"ED8E00",X"FD8F04",X"F98F07",X"F99211",X"FB9519",X"FF9C26",X"EB8C20",X"D07C1C",X"CC802A",X"652904",X"2B0200",X"110400",X"020D11",X"0F2B37",X"123E59",X"3571A3",X"2D76BB",X"1B6ED6",X"0664D5",X"066FEC",X"0776F9",X"0474F2",X"0775E8",X"0069D3",X"137DE3",X"234FA8",X"000020",X"52122A",X"7F1351",X"3F0033",X"0E0011",X"333659",X"113581",X"D5D6EB",X"FBFFFF",X"F3F9F9",X"FAFFF7",X"FCFFF4",X"F9FAF2",X"FFFEFD",X"FFFDFF",X"EDF9FF",X"F6F7E7",X"9997A2",X"0D000E",X"252229",X"0F0004",X"351E0C",X"9A7356",X"D99149",X"F98A2E",X"EC751B",X"E67318",X"E47614",X"FFC886",X"FFFFF0",X"F9FDFC",X"FFFDF7",X"FFFCF9",X"FFFDF9",X"FFFFFA",X"FFFFFA",X"FFFFFB",X"FDFFFA",X"FAFFF9",X"FFFDFE",X"FFFEFD",X"FFFCFB",X"FFFFFF",X"FDFEFF",X"FDFEFF",X"FFFFFA",X"FAF1E8",X"EC7B41",X"F2831A",X"F4792C",X"FF8629",X"F9781A",X"FF7F13",X"FF7C15",X"FF7714",X"FF7B1F",X"F76D00",X"D16A0D",X"FFDFB2",X"FFFFF4",X"FFFDEE",X"FDF7E7",X"F8FFFB",X"F2FFF1",X"FDFDFB",X"FFEDF1",X"E0A583",X"C47B2E",X"C57E48",X"5E2D26",X"110000",X"1A130B",X"060300",X"110D00",X"9C9708",X"F0E82E",X"DEDB10",X"E4DE7C",X"FAF5F1",X"FEFFF5",X"F1FDEF",X"F6F5F3",X"FDF8DA",X"EEB889",X"DB791E",X"F69336",X"FA9744",X"F18E29",X"EE8D2C",X"E79033",X"E79645",X"DF9856",X"C08656",X"885D3A",X"917357",X"F0F7E5",X"F5FFF7",X"F6FFFF",X"F7FFFF",X"FCFFF8",X"FFFFF2",X"FFFFF4",X"FEFDF8",X"EFFFFF",X"FCFFFF",X"FFF9FF",X"FFFBFF",X"FBFFFF",X"F8FFFE",X"FFFBFD",X"FEE7EF",X"B74658",X"860615",X"832933",X"410C1E",X"270D1A",X"000D00",X"062805",X"4F815B",X"7DB983",X"7DC681",X"47884E",X"DBF9E1",X"FAFCFB",X"F6F7F2",X"FFFFFB",X"FFFBFF",X"F9FFFF",X"F6F9FF",X"FFFFFD",X"FDF8F4",X"FDF8F5",X"999B8E",X"000900",X"000A20",X"000E41",X"0D468D",X"2272D3",X"005CCB",X"1572DA",X"1D5EAE",X"000C40",X"0B0425",X"060000",X"9A6641",X"F18C3C",X"F47709",X"FF8813",X"FF8616",X"ED7514",X"F17A26",X"854309",X"4B2A17",X"030504",X"476146",X"7FA870",X"65985D",X"5F995C",X"629A53",X"549E53",X"4F9652",X"5DA364",X"5FA95E",X"4B9A3F",X"64AD51",X"67A154",X"6C9C60",X"5CA64D",X"74B46A",X"74A56E",X"78996A",X"61784C",X"000700",X"000211",X"000027",X"051A53",X"000631",X"01000C",X"9F7660",X"DA8951",X"F88E40",X"F98C37",X"EC8833",X"E39447",X"C28860",X"6A5345",X"000700",X"000800",X"1B1500",X"856113",X"CD9826",X"C3A900",X"DEBF16",X"CAA703",X"CAAB03",X"D3B90C",X"CBB308",X"CFB111",X"D9B320",X"D3A615",X"D1B111",X"CFB90B",X"D2B907",X"C39C00",X"D1A30F",X"C8A418",X"CCB52B",X"D0B252",X"998562",X"010B0A",X"001019",X"4D476B",X"641E5A",X"A23171",X"9B1D67",X"B2237F",X"AD1373",X"B30A6F",X"C20F77",X"C40A77",X"C20375",X"C50076",X"CB017B",X"C6117A",X"BB0375",X"BD1181",X"A42576",X"5A163B",X"000005",X"0C4A49",X"38A1A4",X"00A88D",X"00A489",X"00A48A",X"06AC94",X"09AB94",X"0CA893",X"18AD9A",X"1AAB9A",X"0F9179",X"A2F2E5"),
(X"FAFFE2",X"F1DD7C",X"F4C209",X"E7BF0F",X"E8BD00",X"E7C00D",X"F6CE00",X"EAD200",X"F0D001",X"F7CD19",X"F2BE10",X"FAC612",X"F1C210",X"ECC506",X"EECC08",X"EEC919",X"C7C707",X"FFD016",X"DBB838",X"1D2B00",X"010500",X"12121A",X"001222",X"005D65",X"22CED0",X"1FD6DE",X"0CD0DE",X"10D9E9",X"0CD7E6",X"00C9D3",X"00D3DA",X"06DDE2",X"06D2DD",X"06D6E0",X"00D5DD",X"01D6DC",X"05CED5",X"1FCDD8",X"37C4D6",X"48BCD5",X"4B5A6D",X"00040F",X"090F0D",X"000900",X"27511F",X"78AF6B",X"87BD6F",X"7FAE5E",X"79A75C",X"78B46A",X"62A965",X"77BB80",X"87B688",X"7F987B",X"000500",X"040807",X"110000",X"220000",X"AF671D",X"E88720",X"FF9717",X"F08700",X"FF9F06",X"F79800",X"FF960B",X"F98F07",X"F48D0C",X"F08A0E",X"FF9A24",X"F29327",X"ED9939",X"ECA04A",X"CD916C",X"6A412B",X"0D0000",X"00060A",X"000713",X"000A25",X"00295B",X"0A5398",X"1A6DD5",X"1977E8",X"0C75F2",X"0574F7",X"006EEC",X"0A78EB",X"046FD9",X"0973D9",X"2652AB",X"000020",X"511129",X"A63A78",X"6F2A63",X"0C000F",X"05082B",X"092D79",X"CCCDE2",X"F6FAFF",X"F3F9F9",X"FBFFF8",X"FCFFF4",X"FDFEF6",X"FFFEFD",X"FEF8FC",X"F4FFFF",X"FFFFF1",X"8B8994",X"110012",X"28252C",X"16000B",X"120000",X"280100",X"A25A12",X"E07115",X"F98228",X"F78429",X"E67816",X"FFC987",X"FFFDEE",X"FCFFFF",X"FFFDF7",X"FFFCF9",X"FFFDF9",X"FFFEF9",X"FFFFFA",X"FEFFFA",X"FCFEF9",X"F9FEF8",X"FEFCFD",X"FFFEFD",X"FFFBFA",X"FFFFFF",X"FDFEFF",X"FCFDFF",X"FFFEF9",X"FAF1E8",X"E5743A",X"E97A11",X"EF7427",X"F47518",X"F06F11",X"F97509",X"FD720B",X"FF6F0C",X"FF7A1E",X"FF7609",X"DA7316",X"FFE5B8",X"FFFFF4",X"FFFFF1",X"FCF6E6",X"F8FFFB",X"F7FFF6",X"FFFFFD",X"F4D7DB",X"864B29",X"702700",X"732C00",X"230000",X"130000",X"080100",X"494623",X"AEAA6B",X"DDD849",X"EAE228",X"D7D409",X"FFFA98",X"FFFEFA",X"FBFDF2",X"F8FFF6",X"FFFFFD",X"FFFCDE",X"F2BC8D",X"E17F24",X"FA973A",X"E68330",X"E07D18",X"D27110",X"D67F22",X"A95807",X"762F00",X"5B2100",X"2C0100",X"A28468",X"F8FFED",X"F6FFF8",X"F7FFFF",X"F8FFFF",X"FAFFF6",X"FEFFF1",X"FFFFF4",X"FFFFFA",X"EFFFFF",X"FCFFFF",X"FFF8FF",X"FFFBFF",X"FAFEFF",X"F7FFFD",X"FFFCFE",X"FFE8F0",X"AE3D4F",X"810110",X"520002",X"430E20",X"110004",X"364433",X"769875",X"80B28C",X"5D9963",X"60A964",X"6EAF75",X"CEECD4",X"FEFFFF",X"FFFFFB",X"FFFEFA",X"FFFAFF",X"F4FCFF",X"FBFEFF",X"F6F5F3",X"FFFEFA",X"FFFBF8",X"737568",X"000400",X"0F1A30",X"133B6E",X"2760A7",X"0858B9",X"0163D2",X"0D6AD2",X"2C6DBD",X"243B6F",X"0E0728",X"0D0405",X"2F0000",X"E47F2F",X"FF8214",X"FA7B06",X"FF8717",X"EC7413",X"F67F2B",X"C07E44",X"684734",X"000100",X"000F00",X"729B63",X"619459",X"659F62",X"69A15A",X"57A156",X"68AF6B",X"53995A",X"5DA75C",X"5AA94E",X"59A246",X"6FA95C",X"659559",X"60AA51",X"60A056",X"5E8F58",X"375829",X"000E00",X"000600",X"000312",X"302F5B",X"394E87",X"04133E",X"080413",X"391000",X"D4834B",X"F18739",X"F48732",X"F18D38",X"C8792C",X"310000",X"120000",X"141C07",X"495734",X"878151",X"C8A456",X"E1AC3A",X"BBA100",X"DBBC13",X"DAB713",X"C6A700",X"CFB508",X"CCB409",X"C9AB0B",X"D5AF1C",X"CA9D0C",X"DEBE1E",X"CDB709",X"D7BE0C",X"D7B00D",X"E0B21E",X"E8C438",X"D0B92F",X"705200",X"120000",X"0F1918",X"000710",X"181236",X"6C2662",X"871656",X"81034D",X"8B0058",X"AB1171",X"C0177C",X"B30068",X"B60069",X"D31486",X"CE087F",X"CC027C",X"C9147D",X"C70F81",X"B00474",X"971869",X"350016",X"000005",X"468483",X"319A9D",X"09B398",X"00A88D",X"009F85",X"02A890",X"18BAA3",X"1DB9A4",X"16AB98",X"15A695",X"03856D",X"A6F6E9"),
(X"F8FFE6",X"F1D87E",X"F2C315",X"E6BD0B",X"E3BD02",X"EDBD1B",X"F1C00B",X"E5C30C",X"E4C610",X"EAC602",X"E9BC00",X"F3C404",X"F4CC00",X"F6D106",X"F3CD14",X"EDC808",X"F1CD07",X"F1D12E",X"B69838",X"050300",X"1D140B",X"00140F",X"001B12",X"00080C",X"1D564F",X"4BB8B2",X"30D3D2",X"14D0DB",X"0DD2E3",X"07D4E5",X"10DFEF",X"00C9DB",X"0AD1D8",X"15DAE3",X"09CDD9",X"0CD2DF",X"08D2DE",X"07D3DE",X"00CED4",X"15E4EA",X"1DDCD7",X"009496",X"00424B",X"000B17",X"040002",X"453E2C",X"899B71",X"92BE83",X"6EB164",X"73B164",X"7EB967",X"71AF5A",X"6AA958",X"7AB571",X"70A06E",X"375B37",X"000100",X"090504",X"0E0100",X"583E2D",X"B18A61",X"DB9F59",X"E38E31",X"F69024",X"FB8603",X"FF8F0D",X"FA8D0A",X"FF9710",X"FF9910",X"F6950A",X"E88B00",X"EB8F06",X"FF9C1D",X"F0942D",X"AB5D12",X"813B07",X"4C0C00",X"470D00",X"2E0000",X"210000",X"142431",X"364F6D",X"335C90",X"366BB7",X"2E6EC8",X"2368CF",X"2674E0",X"1C70E0",X"1A68B2",X"09052A",X"560023",X"B9126A",X"CA1274",X"7D0C37",X"1C0000",X"000219",X"DCDCE6",X"FCFFFF",X"FAFFFA",X"F7FDFD",X"F7FAFF",X"FDFBFF",X"FFFDFF",X"FFFEFB",X"FFF4F8",X"EDFFF6",X"78A6DA",X"0053B2",X"2B7AE3",X"003A90",X"000F40",X"000322",X"000313",X"351D1D",X"7D514E",X"9B6A5C",X"956243",X"F0D6C7",X"FDFBFF",X"FFF6FF",X"FEFEFE",X"FDFDFD",X"FDFDFD",X"FEFCFD",X"FFFDFE",X"FFFDFE",X"FDFBFC",X"FCFAFB",X"FFFBFA",X"FFFDFC",X"FDFCFA",X"FDFEFF",X"FAFEFF",X"FCFDFF",X"FFFDF9",X"FDF0E7",X"F9832B",X"EF7D00",X"FD8023",X"ED740B",X"F07D13",X"E77A05",X"EB7D0A",X"EF7F0F",X"E1820E",X"E9871C",X"C87D39",X"F8E2CA",X"F0F6F2",X"FFFFFA",X"FFFCFF",X"FFFBFF",X"FFF7FF",X"FFF7FA",X"A7A5AA",X"070800",X"0B1100",X"040800",X"101000",X"333600",X"B3A20A",X"E3CC40",X"FBE82C",X"F5DF0F",X"EFDB08",X"EED96E",X"FCF8C9",X"F6FFF8",X"FFF2F2",X"FFFEFF",X"FBFFFF",X"EAF7ED",X"AB8875",X"65421A",X"6B532F",X"3F3319",X"3B0409",X"2C0000",X"330000",X"2B0000",X"2C0000",X"3E0B14",X"1E0000",X"C0A0AD",X"FFFBFF",X"FFF9FF",X"FFFBFF",X"FFFAFF",X"FFF9FF",X"FFF9FD",X"FFFBFF",X"FDFDFF",X"FFF8FC",X"FFF9FF",X"FFF6FF",X"FFFAFF",X"FBFCFF",X"FAFEFF",X"FFFEFF",X"FAEEF2",X"675058",X"140000",X"262719",X"000600",X"3F5F4A",X"7AA877",X"7EAF6D",X"5E904B",X"5E934D",X"6BA858",X"619251",X"E1EFD6",X"FFFEFB",X"FDFCF8",X"F5F7F4",X"FFFDFF",X"FBFFFF",X"FEFDFF",X"FFFDFD",X"FFFBF9",X"FFFAFE",X"5D5E72",X"000536",X"293685",X"256ECD",X"1260C4",X"156DD7",X"0567D6",X"0061D0",X"095CC4",X"2564C3",X"0D3B93",X"000315",X"030004",X"704326",X"DA823A",X"F98D28",X"EF8314",X"F98413",X"FD7601",X"F77912",X"AE5B17",X"210000",X"030013",X"2F3E43",X"73966E",X"6FA05F",X"73AB6A",X"4E9B4D",X"5EA360",X"63A064",X"619B5E",X"6BA45F",X"629751",X"679555",X"769D66",X"758966",X"687363",X"000009",X"000019",X"00012A",X"001F5D",X"0A469C",X"1B63CF",X"1A61CB",X"1B4F9A",X"000C2A",X"110000",X"6E3D36",X"DCA297",X"C69181",X"91644D",X"010900",X"040200",X"120200",X"7F670F",X"D7B933",X"CEAB11",X"D0AA0B",X"D5AF0E",X"E3B200",X"E1B717",X"E5C437",X"BFA21A",X"CDAB14",X"D6AF0A",X"D4A801",X"CEA100",X"CAAB03",X"E9BD1C",X"D69F07",X"CE9D14",X"D3B543",X"AA9A4D",X"877B53",X"4E4033",X"000110",X"0D2259",X"06276A",X"000F48",X"001854",X"00154A",X"000432",X"21124B",X"4B3252",X"3C183C",X"57244F",X"743667",X"783266",X"6D2058",X"6B1552",X"B75D9D",X"C14287",X"990B57",X"AB286C",X"5A0C34",X"0A0005",X"001812",X"148D7E",X"0DC0AD",X"0C9585",X"0CA18D",X"09A892",X"029D8B",X"16A496",X"26ACA1",X"1FA99C",X"23B7A7",X"039487",X"A3FBFC"),
(X"FCFFEA",X"ECD379",X"F3C416",X"EDC412",X"ECC60B",X"EFBF1D",X"E8B702",X"E0BE07",X"E4C610",X"EAC602",X"ECBF00",X"EEBF00",X"EFC700",X"F5D005",X"F0CA11",X"E9C404",X"F1CD07",X"EDCD2A",X"755700",X"030100",X"20170E",X"2D4C47",X"204138",X"001317",X"00120B",X"00625C",X"33D6D5",X"20DCE7",X"05CADB",X"0EDBEC",X"00CFDF",X"0BD4E6",X"0AD1D8",X"04C9D2",X"11D5E1",X"0CD2DF",X"02CCD8",X"0AD6E1",X"0EDDE3",X"03D2D8",X"0ECDC8",X"3AD4D6",X"58B2BB",X"14303C",X"050003",X"0D0600",X"1A2C02",X"628E53",X"7ABD70",X"7CBA6D",X"6EA957",X"76B45F",X"7AB968",X"6EA965",X"80B07E",X"88AC88",X"696D6C",X"262221",X"0C0000",X"140000",X"220000",X"9C601A",X"DF8A2D",X"FB9529",X"FF8B08",X"F78604",X"F88B08",X"FC940D",X"F69007",X"F7960B",X"FEA116",X"F79B12",X"F49112",X"E88C25",X"EC9E53",X"DF9965",X"CB8B65",X"8D533B",X"5F2F25",X"290001",X"000310",X"000624",X"00275B",X"063B87",X"2060BA",X"2368CF",X"1D6BD7",X"267AEA",X"1260AA",X"020023",X"5C0629",X"BF1870",X"CF1779",X"9D2C57",X"2D0510",X"060E25",X"D6D6E0",X"FCFFFF",X"F6FDF6",X"F3F9F9",X"FCFFFF",X"FFFDFF",X"FDF8FF",X"FFFEFB",X"FFF9FD",X"ECFFF5",X"72A0D4",X"146BCA",X"2574DD",X"2470C6",X"2C5283",X"324766",X"253646",X"140000",X"1F0000",X"250000",X"350200",X"E1C7B8",X"FFFDFF",X"FFF9FF",X"FDFDFD",X"FDFDFD",X"FCFCFC",X"FEFCFD",X"FFFDFE",X"FEFCFD",X"FDFBFC",X"FBF9FA",X"FFFBFA",X"FFFCFB",X"FCFBF9",X"FDFEFF",X"FAFEFF",X"FCFDFF",X"FFFDF9",X"FDF0E7",X"F9832B",X"F07E00",X"F87B1E",X"FA8118",X"F17E14",X"F58813",X"EA7C09",X"FC8C1C",X"EB8C18",X"E68419",X"C57A36",X"FFEAD2",X"FBFFFD",X"FFFFFA",X"FFFBFF",X"FCF8FF",X"FFF6FF",X"F7EEF1",X"2D2B30",X"000100",X"262C06",X"7F8351",X"A0A05A",X"CBCE5B",X"F7E64E",X"EFD84C",X"EDDA1E",X"F7E111",X"E4D000",X"FDE87D",X"FFFCCD",X"F6FFF8",X"FFFBFB",X"F7F5FA",X"F7FBFF",X"EFFCF2",X"7E5B48",X"1D0000",X"1D0500",X"0B0000",X"2D0000",X"3C0508",X"380104",X"4A1215",X"561D23",X"622F38",X"441A26",X"DBBBC8",X"FFFBFF",X"FFF6FF",X"FFFAFF",X"FFFAFF",X"FFFBFF",X"FFFAFE",X"FEF9FF",X"FAFAFF",X"FFF9FD",X"FFF9FF",X"FFF5FE",X"FFF9FF",X"FBFCFF",X"FAFEFF",X"FFFEFF",X"FBEFF3",X"624B53",X"110000",X"010200",X"46574D",X"80A08B",X"7BA978",X"619250",X"83B570",X"7BB06A",X"5B9848",X"639453",X"DFEDD4",X"FEF9F6",X"FFFEFA",X"FEFFFD",X"FFFCFF",X"F6FBFF",X"FFFEFF",X"FDF7F7",X"FFF9F7",X"FFFDFF",X"636478",X"000233",X"4E5BAA",X"236CCB",X"1462C6",X"0860CA",X"1072E1",X"0466D5",X"1063CB",X"2261C0",X"2351A9",X"011224",X"070208",X"260000",X"C56D25",X"FA8E29",X"EF8314",X"F37E0D",X"FF7B06",X"F67811",X"D78440",X"684438",X"141124",X"000409",X"557850",X"72A362",X"5D9554",X"5DAA5C",X"559A57",X"6EAB6F",X"599356",X"5E9752",X"73A862",X"77A565",X"5B824B",X"344825",X"000500",X"0B0E17",X"000019",X"22315A",X"2F5593",X"205CB2",X"165ECA",X"145BC5",X"3367B2",X"223553",X"0D0000",X"340300",X"82483D",X"632E1E",X"230000",X"000400",X"666457",X"827250",X"C1A951",X"CAAC26",X"CCA90F",X"D7B112",X"D9B312",X"D6A500",X"D3A909",X"C2A114",X"CFB22A",X"C8A60F",X"C8A100",X"EABE17",X"E3B612",X"C4A500",X"E6BA19",X"DAA30B",X"E1B027",X"C5A735",X"78681B",X"1A0E00",X"0B0000",X"181B2A",X"152A61",X"325396",X"1A3972",X"1F3773",X"0A1F54",X"00012F",X"261750",X"4C3353",X"220022",X"2E0026",X"480A3B",X"4F093D",X"41002C",X"3C0023",X"9F4585",X"CE4F94",X"91034F",X"961357",X"4D0027",X"0A0005",X"1C4B45",X"179081",X"00A491",X"0D9686",X"00937F",X"009F89",X"009583",X"069486",X"1AA095",X"149E91",X"15A999",X"009184",X"9AF2F3"),
(X"FAFBFF",X"DBC89D",X"CDB748",X"E6D255",X"D7CA3E",X"E1C243",X"E8CA38",X"E2C931",X"E9CE29",X"EACC12",X"ECCA10",X"E8C60F",X"EDCC0D",X"E6C40B",X"E9C50F",X"E8C300",X"F9C72A",X"CDBC62",X"080C00",X"080000",X"093341",X"1C5B50",X"175957",X"173942",X"001D11",X"000509",X"1C4853",X"4BB8BB",X"31CDCC",X"13C0C7",X"16D6E3",X"01DFEA",X"00D1D6",X"04D5DC",X"01D1DB",X"0ADAE6",X"0BD7E2",X"02CED5",X"0AD7DA",X"07D7D7",X"04D3DD",X"06CCD5",X"20D5E0",X"33C1CF",X"004E5F",X"001021",X"000010",X"080009",X"303636",X"8C9A89",X"9CBC8D",X"73A55E",X"77B761",X"74BA62",X"68AD5C",X"75B86B",X"7BC384",X"70A879",X"2E4E36",X"000400",X"040000",X"100000",X"584026",X"A28563",X"CB8C45",X"DE9340",X"E78B26",X"F28913",X"FC8B0B",X"FF8E0C",X"FF9514",X"FF9616",X"FD8E09",X"F38804",X"FD9613",X"F4910F",X"FD9A22",X"FC9A37",X"DF7D36",X"B65423",X"A35733",X"5F2406",X"190000",X"0B0300",X"000406",X"16293A",X"193155",X"3E5A8A",X"3A4C74",X"000112",X"4B0A2C",X"C91775",X"C60272",X"D21A7A",X"A9054E",X"8D5475",X"FBF1F2",X"FFF9F6",X"FFFFFA",X"FFFEFF",X"FCFAFF",X"FDFBFF",X"FFFEFF",X"FEFEF2",X"FFF9FF",X"D7FFFF",X"559DE7",X"0070DA",X"1478E8",X"0A74E2",X"1774DE",X"1B7FF1",X"106DCD",X"0B4C9E",X"07377F",X"000A40",X"284A65",X"C8ECFA",X"E7FFFF",X"EEFDFF",X"F3FCFF",X"F9FFFF",X"FAFDFF",X"FAF9FF",X"FFFCFF",X"FFF8FF",X"FFF1FF",X"FFF8FF",X"FBFBFD",X"FFFEFF",X"FCFAFB",X"FDFDFF",X"FCFFFF",X"FCFDFF",X"FFFCF8",X"FCEFE6",X"DD996C",X"C38228",X"C97D49",X"C37A47",X"BC7853",X"BA7F55",X"A87148",X"855024",X"8B5D4E",X"714636",X"351508",X"F0E6DD",X"FCFFFD",X"F3F9F9",X"FFFDFF",X"FFF9FF",X"F3FFF3",X"CACF7F",X"6A5E00",X"B29A12",X"DCC52A",X"F6E53D",X"EAE026",X"F9F41C",X"E4D314",X"E9DA0F",X"E3D802",X"EEEB00",X"DFD444",X"FAEDB8",X"FFFBFF",X"F6FDF6",X"FFFEFF",X"FBF7FF",X"FFFBFF",X"F8DAE2",X"A62B3D",X"7A000F",X"910528",X"82002A",X"8B0020",X"9D082E",X"A70D2F",X"AC0928",X"BC0F2D",X"CA1935",X"A90015",X"FF788E",X"FFD5E0",X"FFDCE7",X"FFD2E0",X"FFD4E3",X"FFD6E6",X"FFD3E5",X"FFD6E8",X"FFDDF0",X"FFDBE7",X"FFE6EE",X"FFF5FA",X"FEFCFF",X"F9F8FD",X"FFFDFF",X"FFFEFF",X"F1F3F0",X"43574E",X"000F00",X"5F8959",X"73A373",X"649E64",X"5D9B4E",X"549841",X"7FC272",X"8DC274",X"5E9541",X"668D4C",X"DBE0C9",X"FFFCFD",X"FEFFFA",X"F8FEFA",X"FFFEFF",X"FFFDFF",X"FFF8FB",X"FFFDFD",X"F9FEFA",X"E3FDFE",X"4D7DA3",X"0950A2",X"196ED9",X"0565D6",X"0968D4",X"0D6DD4",X"0263CE",X"0165D5",X"0767DF",X"035DD7",X"1265DD",X"154F8E",X"000329",X"1D111B",X"432314",X"B27E4C",X"F6A147",X"FB8815",X"F77700",X"F97918",X"FA8223",X"C25F1E",X"844639",X"432F3A",X"000600",X"6F9469",X"79A66B",X"63994D",X"6EA250",X"679443",X"6B954D",X"779C69",X"7A967D",X"415147",X"000200",X"050409",X"090C1B",X"021033",X"0F2D69",X"3B6FC3",X"1765C9",X"005FC7",X"0070D7",X"0B6AE2",X"0E63C0",X"2E6EAC",X"000F39",X"000826",X"01000B",X"0A0400",X"39360D",X"654400",X"B9972B",X"E4BF32",X"CBA208",X"E0B818",X"D1B10E",X"C8AF17",X"C7B12A",X"CFAC1E",X"D9B11C",X"CEA307",X"CFA709",X"D3B217",X"CBAE15",X"C5A80E",X"DBBA1D",X"BB9E05",X"D6C144",X"C4B65E",X"9C9159",X"3B3215",X"020202",X"000C2F",X"15326E",X"1850A3",X"1A5CCC",X"125CC7",X"266DC5",X"1259B3",X"1360B8",X"175AB1",X"214EB5",X"053178",X"00165C",X"00094C",X"000340",X"05194C",X"2E3F6B",X"000228",X"000022",X"2D1640",X"441B3D",X"30061A",X"1B0A12",X"000107",X"324E52",X"55988F",X"29937C",X"328C83",X"2E8D85",X"1B897E",X"1C9C8D",X"1BAD9A",X"009C86",X"0BAB91",X"0CAC92",X"058D7F",X"ABF7F7"),
(X"FCFDFF",X"AB986D",X"402A00",X"8E7A00",X"928500",X"C0A122",X"BC9E0C",X"C9B018",X"EED32E",X"E7C90F",X"EFCD13",X"EFCD16",X"E2C102",X"E5C30A",X"EDC913",X"E7C200",X"FFD033",X"96852B",X"000400",X"1A0E10",X"1C4654",X"155449",X"1B5D5B",X"2E5059",X"153327",X"0B1D21",X"000C17",X"005457",X"2FCBCA",X"35E2E9",X"00BECB",X"09E7F2",X"0EDFE4",X"00C7CE",X"0BDBE5",X"07D7E3",X"01CDD8",X"0CD8DF",X"04D1D4",X"0CDCDC",X"10DFE9",X"0ED4DD",X"16CBD6",X"3ECCDA",X"52AFC0",X"2F5A6B",X"040B1B",X"060007",X"000303",X"000C00",X"658556",X"86B871",X"83C36D",X"6AB058",X"6FB463",X"72B568",X"5DA566",X"82BA8B",X"87A78F",X"879188",X"443F39",X"0E0000",X"140000",X"180000",X"5F2000",X"AA5F0C",X"F39732",X"FD941E",X"F07F00",X"FF9513",X"F88B0A",X"FE9313",X"FD8E09",X"F48905",X"FF9B18",X"F99614",X"F5921A",X"F08E2B",X"F08E47",X"EF8D5C",X"E19571",X"B77C5E",X"583821",X"342C21",X"000204",X"000D1E",X"000327",X"000636",X"00062E",X"000314",X"3E001F",X"BB0967",X"D81484",X"D82080",X"AC0851",X"C48BAC",X"FBF1F2",X"FFF9F6",X"FFFFFA",X"FFFEFF",X"FCFAFF",X"FDFBFF",X"FFFEFF",X"FEFEF2",X"FFF7FF",X"CBF3FD",X"2F77C1",X"0068D2",X"0D71E1",X"0B75E3",X"1673DD",X"0E72E4",X"217EDE",X"2F70C2",X"3666AE",X"30598F",X"3F617C",X"97BBC9",X"99B9C4",X"ADBCBF",X"B7C0C5",X"ADB4BA",X"AEB1B8",X"B5B4BC",X"B9B3BF",X"C0B4C2",X"C3B5C4",X"BEADBD",X"EDEDEF",X"FFFDFE",X"FCFAFB",X"FDFDFF",X"FCFFFF",X"FCFDFF",X"FFFEFA",X"FEF1E8",X"8E4A1D",X"7C3B00",X"702400",X"5A1100",X"5C1800",X"541900",X"400900",X"350000",X"220000",X"250000",X"1C0000",X"EBE1D8",X"FCFFFD",X"FBFFFF",X"FFFAFF",X"FFFAFF",X"F1FDF1",X"D8DD8D",X"DFD359",X"F4DC54",X"FBE449",X"E0CF27",X"EBE127",X"E5E008",X"F2E122",X"E8D90E",X"F0E50F",X"E7E400",X"F7EC5C",X"FFF9C4",X"FCF4FF",X"FBFFFB",X"FDFBFC",X"FEFAFF",X"FFFAFF",X"F6D8E0",X"9F2436",X"95142A",X"A81C3F",X"9F1747",X"A7153C",X"A10C32",X"A70D2F",X"B91635",X"B20523",X"B70622",X"B40820",X"BB152B",X"833B46",X"934D58",X"964F5D",X"9A505F",X"994B5B",X"9D5062",X"975264",X"8C4D60",X"9A5E6A",X"724A52",X"BEAFB4",X"FFFEFF",X"FFFEFF",X"FDFBFE",X"FCFAFB",X"F3F5F2",X"70847B",X"729775",X"7AA474",X"77A777",X"659F65",X"70AE61",X"68AC55",X"599C4C",X"6BA052",X"669D49",X"759C5B",X"E5EAD3",X"FFFCFD",X"FDFEF9",X"FBFFFD",X"FAF9FF",X"FFFCFF",X"FFF7FA",X"FFFCFC",X"FAFFFB",X"E9FFFF",X"5888AE",X"135AAC",X"1E73DE",X"0868D9",X"0867D3",X"0767CE",X"0162CD",X"0063D3",X"0464DC",X"0761DB",X"1366DE",X"1F5998",X"162E54",X"070005",X"1D0000",X"75410F",X"F39E44",X"FA8714",X"F77700",X"FB7B1A",X"F27A1B",X"E3803F",X"A26457",X"0D0004",X"000600",X"0C3106",X"6D9A5F",X"699F53",X"689C4A",X"7BA857",X"749E56",X"456A37",X"132F16",X"000600",X"000503",X"06050A",X"191C2B",X"101E41",X"4765A1",X"3064B8",X"1462C6",X"056AD2",X"0063CA",X"005FD7",X"085DBA",X"2262A0",X"385D87",X"00011F",X"181422",X"332D1D",X"88855C",X"D5B467",X"C8A63A",X"C49F12",X"CFA60C",X"E2BA1A",X"CBAB08",X"BEA50D",X"C7B12A",X"DFBC2E",X"CFA712",X"DCB115",X"D7AF11",X"C7A60B",X"CFB219",X"EFD238",X"C7A609",X"E0C32A",X"B29D20",X"978931",X"130800",X"0A0100",X"191919",X"1E2C4F",X"3A5793",X"2B63B6",X"1C5ECE",X"1E68D3",X"1960B8",X"165DB7",X"1562BA",X"2265BC",X"2D5AC1",X"335FA6",X"375CA2",X"385396",X"354986",X"425689",X"2F406C",X"1A264C",X"0D1337",X"0B001E",X"1C0015",X"1D0007",X"0B0002",X"000107",X"001519",X"0B4E45",X"005B44",X"005A51",X"207F77",X"158378",X"058576",X"089A87",X"0CA892",X"009F85",X"0EAE94",X"00887A",X"A8F4F4"),
(X"FFF3FF",X"978E93",X"000700",X"000300",X"000402",X"030004",X"14110C",X"281B13",X"573C1F",X"AF9155",X"F0CF4A",X"EED00E",X"EBCC00",X"E4C300",X"EDC605",X"F3C321",X"EEC23B",X"534514",X"040809",X"0D271E",X"0C5B55",X"045F5A",X"106464",X"00575E",X"235E64",X"003D3C",X"001919",X"000007",X"223A3C",X"46AEA5",X"35DAD4",X"14C5CB",X"12DBE3",X"00D1D8",X"00D3DC",X"00D7E1",X"02D8E3",X"04D9E1",X"02D7DB",X"04DCDB",X"01D1DD",X"00CFDC",X"10E6F1",X"00DCE4",X"01DADF",X"1CD9DF",X"1CAEBB",X"00465A",X"000D10",X"0C1F26",X"000007",X"4B5453",X"6E8B75",X"7DAD7B",X"89BA6B",X"86AF51",X"6CB367",X"6CAF5F",X"7DBB66",X"88C26D",X"6FA559",X"649158",X"648363",X"000C00",X"000608",X"030100",X"674E2F",X"AF804A",X"DA964D",X"ED9438",X"F98F22",X"FC850F",X"F98E00",X"F68800",X"FF9209",X"FA8F03",X"F69200",X"F29500",X"F29901",X"F09802",X"FF9417",X"FF9620",X"E08115",X"F29E3E",X"AE6719",X"5A2100",X"270000",X"190000",X"250905",X"140000",X"1E0113",X"A52465",X"D80A79",X"E60F90",X"CB097B",X"DF79BA",X"FFEDFF",X"FFF5FF",X"FFFDFB",X"FFFDFA",X"FDFCFF",X"FDFEFF",X"FEFFFD",X"FDFFF2",X"FFF8FF",X"CFE8FC",X"0C65B7",X"0B70E2",X"0075D7",X"0F6ADD",X"0772E6",X"0473F8",X"0074DE",X"016ED7",X"157EE9",X"1074E3",X"156FDF",X"095BC9",X"0148B0",X"003596",X"002A90",X"001675",X"000959",X"000340",X"00052C",X"00061B",X"000A0F",X"000805",X"DCE1E7",X"FAFBFF",X"FEFCFD",X"FFFDFE",X"FEFEFF",X"FCFCFE",X"FFFEFB",X"FBF4EE",X"2F304F",X"030700",X"0A0100",X"0D0300",X"0F0300",X"0B0300",X"0C0500",X"100B00",X"453800",X"574F00",X"615900",X"F9F3B5",X"FFFCF3",X"F9FBFF",X"FDFBEF",X"FFFDCF",X"FFF66B",X"E1D310",X"EFDF06",X"EDD908",X"F1DE05",X"F5DC03",X"FFD90F",X"F7C600",X"EDDD00",X"E8DA08",X"E6E028",X"DDD66C",X"F3F1B8",X"FFFCFF",X"FFFFFF",X"F9FCF5",X"FDFEF6",X"FFFCFF",X"FFFAF8",X"F7CCC6",X"A80108",X"B71223",X"C30921",X"BD0424",X"C00A23",X"C00925",X"BD0423",X"C70528",X"CC052E",X"C10027",X"CD0E39",X"B00023",X"C8071A",X"BD0215",X"B00010",X"B6091D",X"A80218",X"9F061A",X"950B1A",X"870813",X"591E20",X"1A0000",X"A19E99",X"FBFFFF",X"F4F2F5",X"FFFAFF",X"FFFFFD",X"EEFBF2",X"8AA584",X"76B56F",X"689D4F",X"72A55A",X"64A255",X"71B15D",X"55A250",X"5EA964",X"5A9F4E",X"61A751",X"6C9C5E",X"DCEBD6",X"FBFBFD",X"F7FDF9",X"FBFFFD",X"FFFBFF",X"FFFDFD",X"FFFAF8",X"FFFAFF",X"F9FDFE",X"E7FFFF",X"568DC5",X"085AC6",X"096FEB",X"0166D8",X"0066D4",X"0064D1",X"0066D9",X"0067E0",X"0168E1",X"0D67D7",X"0B5DC3",X"1E60D0",X"2F58A8",X"161E43",X"0A0002",X"513834",X"986D5A",X"E7905A",X"F7771E",X"F08924",X"FA841A",X"EF740A",X"DD751C",X"803402",X"491A10",X"060004",X"536D6C",X"93B582",X"769569",X"62795C",X"2A352D",X"030004",X"1A0000",X"491800",X"6C2E00",X"5E310A",X"270E00",X"060D05",X"2A516E",X"1B5C9E",X"1263BF",X"0961C5",X"065FC3",X"115BC4",X"0C67D0",X"0467CF",X"196DCF",X"063881",X"000829",X"090700",X"6E673B",X"C4A241",X"CFB018",X"CCAE00",X"CDA90B",X"D4AF44",X"E8CD80",X"B6A86B",X"686232",X"505443",X"9A9865",X"BCAF47",X"D0B21E",X"D3A905",X"C79E06",X"C3A628",X"C9B44B",X"A49B62",X"453F1F",X"080000",X"0F0009",X"14000E",X"05001A",X"466294",X"306DAE",X"0061B6",X"035CD4",X"0967D9",X"0059B4",X"0061C7",X"0555C6",X"024EBE",X"085DD2",X"0564D8",X"126BDF",X"196DDF",X"196BD7",X"267CDF",X"055CB9",X"0A5EB4",X"0253A5",X"0D48AE",X"00297B",X"002A66",X"002960",X"001F5D",X"000442",X"000734",X"000119",X"010B17",X"060C1C",X"000C1B",X"044446",X"1C9586",X"069E85",X"008F76",X"1F9C8A",X"00876A",X"A6F2E5"),
(X"FFF6FF",X"A49BA0",X"000700",X"212821",X"000402",X"0A050B",X"030000",X"0E0100",X"1A0000",X"301200",X"D3B22D",X"EED00E",X"EACB00",X"EAC900",X"E2BB00",X"FFD230",X"CEA21B",X"150700",X"000102",X"1D372E",X"1A6963",X"06615C",X"0B5F5F",X"0F666D",X"215C62",X"115554",X"0A3232",X"0C0C14",X"00090B",X"00433A",X"23C8C2",X"2EDFE5",X"00C7CF",X"0CDDE4",X"03DCE5",X"00DAE4",X"00CDD8",X"00CED6",X"0FE4E8",X"01D9D8",X"0CDCE8",X"00CBD8",X"03D9E4",X"00DBE3",X"06DFE4",X"14D1D7",X"39CBD8",X"3EADC1",X"41676A",X"000F16",X"000007",X"000403",X"001100",X"477745",X"89BA6B",X"89B254",X"74BB6F",X"61A454",X"6FAD58",X"79B35E",X"7FB569",X"7EAB72",X"9FBE9E",X"657A69",X"000305",X"070500",X"1A0100",X"340500",X"955108",X"DC8327",X"FF9F32",X"FF8913",X"FD9204",X"FB8D02",X"FE9007",X"FD9206",X"F99501",X"F39600",X"EE9500",X"EB9300",X"F38508",X"FF9620",X"EE8F23",X"E69232",X"E9A254",X"CF9661",X"A57B62",X"5A3C32",X"140000",X"22050A",X"1C0011",X"8A094A",X"E21483",X"EF1899",X"BF006F",X"DF79BA",X"FFEEFF",X"FFF6FF",X"FFFDFB",X"FFFDFA",X"FDFCFF",X"FEFFFF",X"FEFFFD",X"FDFFF2",X"FFF8FF",X"C8E1F5",X"0760B2",X"1A7FF1",X"0379DB",X"0A65D8",X"036EE2",X"0776FB",X"067BE5",X"0C79E2",X"026BD6",X"1074E3",X"1670E0",X"1C6EDC",X"2C73DB",X"346ECF",X"3F69CF",X"456DCC",X"3C61B1",X"365895",X"3B5B82",X"324E63",X"274045",X"2D4643",X"DADFE5",X"FBFCFF",X"FFFEFF",X"FFFEFF",X"FEFEFF",X"FDFDFF",X"FFFEFB",X"F9F2EC",X"303150",X"1F2300",X"4C4324",X"5E5421",X"6E623C",X"81794B",X"A09965",X"B4AF6D",X"D7CA62",X"DAD263",X"D5CD68",X"FFFFC1",X"FFFEF5",X"F9FBFF",X"FFFFF4",X"FFF7C9",X"E3D045",X"E9DB18",X"F4E40B",X"F0DC0B",X"E6D300",X"F4DB02",X"F3CC02",X"FFDD14",X"EDDD00",X"EBDD0B",X"EBE52D",X"CFC85E",X"FFFEC5",X"FFFDFF",X"FFFFFF",X"F7FAF3",X"FBFCF4",X"FFFCFF",X"FFFCFA",X"F4C9C3",X"A30003",X"C11C2D",X"C0061E",X"BC0323",X"BC061F",X"C10A26",X"C20928",X"BC001D",X"D00932",X"C30029",X"BE002A",X"C20C35",X"CD0C1F",X"C70C1F",X"C10E21",X"C6192D",X"B91329",X"B0172B",X"A21827",X"890A15",X"5E2325",X"160000",X"94918C",X"FAFFFE",X"FEFCFF",X"FFFCFF",X"FEFEFC",X"EDFAF1",X"90AB8A",X"56954F",X"6CA153",X"689B50",X"5A984B",X"6DAD59",X"529F4D",X"64AF6A",X"66AB5A",X"599F49",X"5E8E50",X"D1E0CB",X"FFFFFF",X"F7FDF9",X"F9FFFB",X"FFFDFF",X"FFFDFD",X"FFFDFB",X"FFFAFF",X"F8FCFD",X"E4FFFF",X"568DC5",X"0355C1",X"0167E3",X"0368DA",X"0064D2",X"0064D1",X"0472E5",X"006CE5",X"0061DA",X"0E68D8",X"1163C9",X"1658C8",X"3059A9",X"2A3257",X"54454C",X"381F1B",X"2B0000",X"CB743E",X"FE7E25",X"FA932E",X"FF9127",X"F0750B",X"EA8229",X"C37745",X"56271D",X"201A1E",X"0D2726",X"577946",X"304F23",X"000A00",X"000400",X"030004",X"1A0000",X"956444",X"CF9158",X"B68962",X"4A3113",X"000400",X"00102D",X"2162A4",X"0D5EBA",X"0159BD",X"0B64C8",X"1660C9",X"035EC7",X"0669D1",X"0F63C5",X"2F61AA",X"071637",X"030100",X"1F1800",X"BB9938",X"D7B820",X"DEC006",X"DEBA1C",X"B59025",X"A98E41",X"5E5013",X"0F0900",X"000300",X"0D0B00",X"978A22",X"D2B420",X"C89E00",X"D5AC14",X"D9BC3E",X"8D780F",X"0D0400",X"0F0900",X"2A1E1E",X"573E51",X"40223A",X"221737",X"173365",X"2E6BAC",X"056BC0",X"0861D9",X"0563D5",X"006AC5",X"0568CE",X"0E5ECF",X"0A56C6",X"075CD1",X"005DD1",X"0057CB",X"085CCE",X"0E60CC",X"156BCE",X"1B72CF",X"0D61B7",X"1667B9",X"1E59BF",X"265DAF",X"2A609C",X"2A5D94",X"325896",X"283A78",X"141F4C",X"27334B",X"000713",X"0B1121",X"000413",X"08484A",X"259E8F",X"029A81",X"08987F",X"25A290",X"00896C",X"A6F2E5"),
(X"EBFFF5",X"87D6C3",X"119F87",X"1D9D8E",X"028D78",X"109077",X"0B9272",X"047257",X"0B2518",X"000300",X"867327",X"F3D040",X"F3CB14",X"E0BA00",X"E9C710",X"EFC83F",X"84774B",X"010204",X"06191F",X"005051",X"0F644F",X"005D62",X"00554D",X"007262",X"006768",X"09585D",X"175B5C",X"00362E",X"001B14",X"00080F",X"063138",X"57B2B3",X"37D1D3",X"19C5C5",X"0DCFD1",X"0EDDE3",X"02D2DE",X"00CAD9",X"0AD5E4",X"08D6E3",X"08D2DC",X"08DEE6",X"00DFE5",X"00D7E0",X"0CD7E6",X"0FCEE0",X"0FD0DF",X"1AE0EB",X"26CCD8",X"0FA5A6",X"00625C",X"001612",X"000A0C",X"0D0405",X"4B5443",X"8EAD8B",X"8AAD77",X"92B87B",X"80AF69",X"74AF5F",X"6FB35C",X"71B65D",X"79B460",X"8EC371",X"779E72",X"3D5F3E",X"000D00",X"000702",X"030E08",X"474225",X"917335",X"CE9E49",X"E99439",X"EC902D",X"EF8B19",X"FB9212",X"FF950B",X"FF940A",X"FF9411",X"FF981B",X"FA9000",X"FA8B00",X"FF8C04",X"FC8000",X"FF8B0A",X"F98C13",X"F59E2D",X"E7A036",X"AF7047",X"220A00",X"110000",X"98104E",X"D91C7A",X"E61283",X"D70069",X"DD87B4",X"FFF0FF",X"FFF7FF",X"FFFDFF",X"FFFEF9",X"FDFEF8",X"FEFFFB",X"FFFFFD",X"FEFDFB",X"FDFEFF",X"B8D9F8",X"0A5DC5",X"187BF3",X"027CE1",X"0A6EE8",X"0070E7",X"0070EC",X"016BDB",X"097CE7",X"0073DA",X"0C7FEA",X"0A77EC",X"056CE3",X"1076E2",X"0A76D8",X"006ADD",X"0A75E7",X"0973E3",X"0D73E1",X"1A7CE7",X"1676DD",X"0F6CD3",X"1975DA",X"D6E2EE",X"FAFEFF",X"FFFEFF",X"FFFDFC",X"FEFCFD",X"FDFDFF",X"FFFFFF",X"F2F1EF",X"1E192D",X"767920",X"DFD854",X"E3D824",X"EEDF2E",X"F3E32E",X"F4E324",X"FEEC1C",X"EEEA05",X"F6E90E",X"F1E53B",X"FAF6AC",X"FBFBFD",X"FFFCF9",X"FFFEB1",X"EBEF5C",X"EADA0B",X"F0E207",X"F0E011",X"E7D712",X"F6EC19",X"EAE510",X"DED70D",X"E5E00B",X"F0DF15",X"FBE947",X"C1AF59",X"E4DAB7",X"FFFAFF",X"FCFDFF",X"FCFDFF",X"FEFCFF",X"FCFDFF",X"FEF9FF",X"FFFDFF",X"F5C7CA",X"B40008",X"CB1C3D",X"CD0023",X"CF0026",X"C70528",X"BC001D",X"C80428",X"C60024",X"C90125",X"C60323",X"B90019",X"B5051A",X"B51133",X"A30E2B",X"95172D",X"8B253A",X"691F2E",X"390B0E",X"230F06",X"191400",X"101000",X"0B1300",X"96A392",X"FAFFFA",X"FFFDFF",X"FFFDFF",X"FCFEFB",X"EDFAF0",X"90AC7C",X"4D9F4A",X"69A84F",X"6CA153",X"609E51",X"6CA254",X"66A658",X"649C5D",X"61A05A",X"5A9A50",X"68945F",X"D0DCD0",X"FEFFFF",X"F6FFFC",X"F5FAF4",X"FFFAFF",X"F9FEF8",X"FFFEFA",X"FFF9FF",X"FFFBFF",X"EDFAFF",X"6588C8",X"134FC7",X"1265DF",X"1564DB",X"0A5ED0",X"0660D0",X"1372E6",X"0B6CDD",X"035DBE",X"1968AB",X"246B97",X"2B4786",X"00173D",X"0E1B14",X"3F2902",X"250D00",X"070002",X"5B3B2E",X"D2854D",X"D18226",X"FB983A",X"ED7C14",X"F6861A",X"EF7E20",X"BE551B",X"5F1B08",X"200308",X"1B0627",X"17000B",X"1C0000",X"320100",X"844404",X"D37E2D",X"F88C32",X"F4791B",X"FF7F34",X"DE7136",X"3B0000",X"1F0C12",X"102854",X"3069B6",X"0957BC",X"0F66DA",X"0A53B9",X"0C62CF",X"0062D7",X"0666DF",X"1562CE",X"2352A0",X"000D37",X"000211",X"767758",X"ACAF78",X"AAAF6C",X"797C4F",X"141613",X"00021F",X"000125",X"001133",X"140E56",X"05002D",X"040000",X"968C51",X"D0C166",X"B1A456",X"7C7757",X"01040B",X"3B1842",X"59084A",X"860258",X"B32579",X"912966",X"2F002B",X"05002A",X"2C3669",X"246EAD",X"1358BD",X"0253BE",X"096AC9",X"0862D2",X"0E5BD1",X"156CD3",X"0062C1",X"0864CB",X"065DC7",X"0E60D0",X"0D5ED1",X"075DCE",X"1A71E2",X"0056C7",X"0C5ECE",X"1A68E4",X"005CC9",X"0266C8",X"0663C3",X"1363C4",X"2D70C7",X"2D5DA5",X"24437C",X"082E31",X"002A30",X"004142",X"25948B",X"009883",X"00A588",X"16BDA1",X"11A990",X"079587",X"ACFCFD"),
(X"F0FFFA",X"77C6B3",X"18A68E",X"3CBCAD",X"2DB8A3",X"36B69D",X"31B898",X"40AE93",X"304A3D",X"080B00",X"5E4B00",X"E8C535",X"F2CA13",X"ECC600",X"EAC811",X"E3BC33",X"2A1D00",X"000002",X"182B31",X"025253",X"055A45",X"04676C",X"025F57",X"007767",X"006263",X"1B6A6F",X"125657",X"1A5B53",X"053029",X"000D14",X"00131A",X"003E3F",X"26C0C2",X"2FDBDB",X"0DCFD1",X"02D1D7",X"11E1ED",X"07D2E1",X"01CCDB",X"02D0DD",X"08D2DC",X"00D1D9",X"00DCE2",X"06E3EC",X"01CCDB",X"11D0E2",X"16D7E6",X"0DD3DE",X"2AD0DC",X"46DCDD",X"43B4AE",X"2F6A66",X"00080A",X"070000",X"000800",X"183715",X"567943",X"7EA467",X"90BF79",X"77B262",X"64A851",X"75BA61",X"72AD59",X"689D4B",X"83AA7E",X"97B998",X"718C7B",X"253A35",X"000400",X"070200",X"1C0000",X"683800",X"C67116",X"ED912E",X"FB9725",X"FA9111",X"F18700",X"F48900",X"FB8C09",X"FD8B0E",X"FF9505",X"FE8F02",X"FF960E",X"FF8F0B",X"FF8A09",X"FF9219",X"E99221",X"E9A238",X"C08158",X"361E06",X"1B010A",X"9C1452",X"CE116F",X"E81485",X"DB026D",X"D57FAC",X"FFF1FF",X"FFF8FF",X"FFFDFF",X"FFFEF9",X"FDFEF8",X"FEFFFB",X"FFFFFD",X"FEFDFB",X"FCFDFF",X"BFE0FF",X"1164CC",X"1679F1",X"037DE2",X"0F73ED",X"0477EE",X"006FEB",X"0670E0",X"0477E2",X"0075DC",X"0376E1",X"0E7BF0",X"0062D9",X"0A70DC",X"0773D5",X"1785F8",X"0D78EA",X"0973E3",X"0B71DF",X"0A6CD7",X"0E6ED5",X"126FD6",X"0F6BD0",X"D7E3EF",X"F9FDFF",X"FFFDFF",X"FFFBFA",X"FEFCFD",X"FDFDFF",X"FFFFFF",X"F2F1EF",X"0C071B",X"767920",X"F6EF6B",X"EFE430",X"EBDC2B",X"EEDE29",X"F1E021",X"F5E313",X"E5E100",X"EADD02",X"E7DB31",X"FFFFB7",X"FFFFFF",X"FFFEFB",X"EBE89B",X"DADE4B",X"F5E516",X"F0E207",X"EEDE0F",X"E8D813",X"ECE20F",X"E2DD08",X"EAE319",X"EAE510",X"F3E218",X"D1BF1D",X"B4A24C",X"FFFFDD",X"FFF9FF",X"FDFEFF",X"FCFDFF",X"FDFBFE",X"FEFFFF",X"FDF8FF",X"FFFDFF",X"F2C4C7",X"B10005",X"C41536",X"C8001E",X"CC0023",X"C40225",X"C20023",X"C70327",X"CE082C",X"CA0226",X"CC0929",X"CB102B",X"B9091E",X"B30F31",X"9B0623",X"810319",X"6E081D",X"631928",X"290000",X"0F0000",X"060100",X"303014",X"596149",X"BAC7B6",X"F8FFF8",X"FCF7FB",X"FFFCFE",X"FEFFFD",X"EFFCF2",X"89A575",X"4EA04B",X"5E9D44",X"6DA254",X"69A75A",X"70A658",X"5E9E50",X"659D5E",X"609F59",X"6BAB61",X"709C67",X"CDD9CD",X"FEFFFF",X"F6FFFC",X"F9FEF8",X"FFFAFF",X"F8FDF7",X"FFFFFB",X"FFF9FF",X"FFFDFF",X"ECF9FF",X"6487C7",X"124EC6",X"1568E2",X"0B5AD1",X"0C60D2",X"0761D1",X"0564D8",X"096ADB",X"126CCD",X"105FA2",X"004470",X"000A49",X"00143A",X"000500",X"69532C",X"5E462E",X"090004",X"190000",X"AD6028",X"EC9D41",X"D67315",X"FF8F27",X"F6861A",X"FF9638",X"E2793F",X"B6725F",X"46292E",X"725D7E",X"110005",X"633F33",X"B4835A",X"CD8D4D",X"FCA756",X"F98D33",X"E86D0F",X"F36F24",X"EF8247",X"8F4E30",X"17040A",X"000632",X"104996",X"1E6CD1",X"085FD3",X"0D56BC",X"1167D4",X"0C6FE4",X"005DD6",X"115ECA",X"3160AE",X"162953",X"00000E",X"070800",X"363902",X"252A00",X"040700",X"000100",X"29304D",X"37476B",X"405779",X"2E2870",X"211B49",X"0B0602",X"544A0F",X"96872C",X"403300",X"070200",X"000007",X"58355F",X"914082",X"9E1A70",X"9E1064",X"912966",X"481744",X"000025",X"000437",X"075190",X"1E63C8",X"0C5DC8",X"0566C5",X"1973E3",X"0956CC",X"136AD1",X"0774D3",X"005CC3",X"085FC9",X"0E60D0",X"095ACD",X"0258C9",X"075ECF",X"0D63D4",X"1567D7",X"1B69E5",X"0059C6",X"0A6ED0",X"0562C2",X"0D5DBE",X"1D60B7",X"1F4F97",X"001D56",X"000B0E",X"0C373D",X"327677",X"1E8D84",X"17B09B",X"00A88B",X"00A68A",X"1BB39A",X"018F81",X"A4F4F5"),
(X"FDFEF6",X"7BD2C2",X"00AF9A",X"16BAA1",X"00B390",X"11BD97",X"0ABEA3",X"27BAB0",X"3B898B",X"000E07",X"090400",X"CBA753",X"F4CB23",X"E1BF06",X"F5D751",X"9F8524",X"000205",X"050700",X"0F3E38",X"186054",X"125A57",X"134C55",X"004E64",X"0A635F",X"005C4F",X"04655E",X"00585D",X"17616E",X"16545F",X"06393C",X"001414",X"000206",X"0D3942",X"5CB1B4",X"46D7D4",X"0BCAC5",X"01D3D4",X"06D9E2",X"0BD6E5",X"03CADD",X"01D1D5",X"0ED9E0",X"0ED4DF",X"08D1DB",X"00CED6",X"05DAE0",X"03D8DE",X"01D2D7",X"00DAE9",X"00CAD5",X"18D7E1",X"2EDAE4",X"0FA1AE",X"004E5B",X"000E15",X"00080A",X"000200",X"2C3425",X"7E926F",X"9ABF89",X"7EB26A",X"6BA85A",X"78B768",X"77B165",X"6BB465",X"67A655",X"89BE6E",X"82B06F",X"638E61",X"1D3D26",X"000500",X"080806",X"030100",X"52422B",X"9A744D",X"CF9556",X"E49A43",X"F19A30",X"F6931C",X"F68D0E",X"FF9E0F",X"F39406",X"F4970B",X"F39406",X"F79003",X"FF960D",X"F88904",X"FF9113",X"EC9F59",X"6C4019",X"120000",X"92135A",X"D5167D",X"F01D88",X"DB005E",X"EB85AD",X"FCF8F7",X"FEFCFF",X"FEFFFF",X"FDFEFF",X"FDFFFE",X"FFFFFF",X"FFFEFF",X"FFFAFF",X"FCFFF6",X"C4E0F6",X"1C42A7",X"2472D6",X"2774CC",X"1271DB",X"1D75DF",X"1477D5",X"0C69E2",X"0773E2",X"0065C9",X"107AE0",X"0A6DE4",X"1573ED",X"016BDB",X"0583EA",X"0674E5",X"006BDC",X"016CDE",X"0671E3",X"0771E1",X"0973E3",X"0971E2",X"0169DA",X"D5E5F5",X"F5FCFF",X"FEFCFF",X"FFFCF9",X"FFFDFC",X"FDFDFD",X"FEFFFF",X"F2F3F5",X"1D0C2E",X"6E6603",X"F1E539",X"F7EB03",X"F0DE02",X"EEDA0A",X"F3DC10",X"F3DC04",X"F4E119",X"FBD906",X"EBD426",X"FBFFAE",X"EEFAEC",X"FEF2E2",X"E0CC91",X"D0CA6C",X"E5DA70",X"DAD168",X"D7CF6D",X"DBD269",X"D7CE59",X"DBCF6D",X"D8CD74",X"D0CD5A",X"E1E787",X"9B986B",X"E8E3DD",X"F9F9F9",X"FBFFF6",X"FBFFFD",X"FBFBF9",X"FFFAF8",X"FFFFF0",X"FFF9FF",X"F9FFF2",X"E8CDC2",X"A30000",X"B1273E",X"B30F27",X"B7132C",X"AC142B",X"AB1832",X"9B152E",X"90162F",X"841A31",X"6F1A2D",X"61232E",X"4D1E24",X"2A1011",X"231411",X"0A0702",X"000400",X"4A5A57",X"5F796E",X"6C9279",X"679771",X"68A770",X"6E9D71",X"ABC3AB",X"FEFFFA",X"FFFEFF",X"FFFDFE",X"F8FDF7",X"F3FDF4",X"8F9F78",X"54A556",X"69A859",X"629955",X"5EA059",X"7AAF5F",X"5E9A44",X"6C9C50",X"7CA16D",X"739A61",X"445D36",X"C0C0BE",X"FDFAFF",X"F7FFFF",X"FCFFFB",X"FFFBFF",X"F7FFFB",X"FEFFFB",X"FFFAFF",X"FEFFFF",X"E4FCFC",X"5A8CC1",X"0453BC",X"0A70D5",X"0063D2",X"0063CB",X"0962C6",X"115CC1",X"215CBA",X"2A529A",X"1C3259",X"111B25",X"271C22",X"040700",X"727800",X"E6E442",X"BAB22B",X"2A2600",X"0B0C00",X"000306",X"C28767",X"F79959",X"F17A2A",X"FF8F44",X"F1832C",X"EF8112",X"E97E16",X"C7651A",X"B66D0E",X"DA812F",X"EC7D38",X"FF853B",X"F4771B",X"E97005",X"F98315",X"F17C12",X"F68609",X"EC8423",X"E28C51",X"652D12",X"0D0000",X"081F3E",X"205599",X"165CBE",X"076AE2",X"0053C0",X"2476DA",X"0D66CE",X"0167D5",X"0161C7",X"2469B4",X"001C4F",X"000017",X"000038",X"00004D",X"001F6B",X"104799",X"195DC2",X"1260CD",X"1F75DC",X"0962C6",X"0D4A9B",X"001C4F",X"00071E",X"00050D",X"07000E",X"4F0B3C",X"8E1C64",X"B10567",X"BE0B73",X"C60578",X"D90985",X"C20070",X"B61D77",X"6E1C4D",X"110007",X"120C30",X"315299",X"1961B6",X"0B5EBE",X"196CE4",X"005AD3",X"0061C5",X"0D71CF",X"0562CC",X"0A62D0",X"095DCD",X"065CCB",X"025CCA",X"0059C1",X"1470D7",X"1A71D8",X"0655BC",X"0B69CD",X"065EC0",X"1955B5",X"4573BE",X"2B5480",X"01172E",X"0A0615",X"002626",X"15726A",X"37BEAD",X"049F8D",X"12AA9B",X"0FA292",X"0FA290",X"15AE99",X"029680",X"A7FCF5"),
(X"FCFDF5",X"80D7C7",X"03B39E",X"1DC1A8",X"0EC29F",X"0DB993",X"04B89D",X"2ABDB3",X"3F8D8F",X"00120B",X"080300",X"9D7925",X"FED52D",X"EDCB12",X"D7B933",X"5D4300",X"000205",X"1D1F12",X"1B4A44",X"125A4E",X"0D5552",X"175059",X"0A5C72",X"035C58",X"035F52",X"006059",X"0A656A",X"06505D",X"25636E",X"1C4F52",X"102E2E",X"0B1014",X"000C15",X"004043",X"2CBDBA",X"26E5E0",X"04D6D7",X"09DCE5",X"04CFDE",X"0FD6E9",X"00CFD3",X"03CED5",X"08CED9",X"0BD4DE",X"0CDBE3",X"05DAE0",X"01D6DC",X"02D3D8",X"00DCEB",X"05D8E3",X"16D5DF",X"19C5CF",X"3ED0DD",X"58C0CD",X"54858C",X"000305",X"020703",X"000500",X"000E00",X"537842",X"79AD65",X"7FBC6E",X"6DAC5D",X"77B165",X"6BB465",X"7AB968",X"77AC5C",X"77A564",X"86B184",X"85A58E",X"64736C",X"363634",X"19170A",X"160600",X"1F0000",X"682E00",X"AE640D",X"D88117",X"F18E17",X"FF9E1F",X"FA9708",X"EE8F01",X"F79A0E",X"F39406",X"FF9B0E",X"FF930A",X"FB8C07",X"F78709",X"E79A54",X"7D512A",X"110000",X"96175E",X"CE0F76",X"EC1984",X"D9005C",X"F08AB2",X"FCF8F7",X"FEFCFF",X"FEFFFF",X"FDFEFF",X"FDFFFE",X"FFFFFF",X"FFFEFF",X"FFFAFF",X"FCFFF6",X"B1CDE3",X"001378",X"1967CB",X"2C79D1",X"1170DA",X"1D75DF",X"187BD9",X"0C69E2",X"0571E0",X"0272D6",X"0872D8",X"096CE3",X"0F6DE7",X"0069D9",X"0381E8",X"0371E2",X"0977E8",X"036EE0",X"006BDD",X"0C76E6",X"0771E1",X"0169DA",X"0A72E3",X"D6E6F6",X"F6FDFF",X"FFFDFF",X"FFFEFB",X"FFFEFD",X"FDFDFD",X"FEFFFF",X"F3F4F6",X"211032",X"7D7512",X"F1E539",X"EBDF00",X"F7E509",X"F4E010",X"F2DB0F",X"FFEA12",X"F2DF17",X"FBD906",X"F2DB2D",X"F9FFAC",X"F5FFF3",X"FFF9E9",X"F6E2A7",X"E9E385",X"F1E67C",X"EBE279",X"F5ED8B",X"EBE279",X"F4EB76",X"F4E886",X"EFE48B",X"EDEA77",X"E3E989",X"F9F6C9",X"FFFCF6",X"FFFFFF",X"F9FFF4",X"F4FAF6",X"FFFFFD",X"FFFDFB",X"FFFDEE",X"FFFCFF",X"F8FFF1",X"EBD0C5",X"9F0000",X"B1273E",X"B00C24",X"B20E27",X"AD152C",X"900017",X"8C061F",X"7F051E",X"70061D",X"540012",X"390006",X"200000",X"140000",X"0B0000",X"080500",X"2B342F",X"95A5A2",X"809A8F",X"769C83",X"80B08A",X"609F68",X"639266",X"A4BCA4",X"FEFFFA",X"FDF9FA",X"FEFCFD",X"FAFFF9",X"F1FBF2",X"94A47D",X"4C9D4E",X"65A455",X"679E5A",X"5EA059",X"659A4A",X"64A04A",X"73A357",X"81A672",X"50773E",X"000C00",X"A7A7A5",X"FFFDFF",X"F9FFFF",X"FAFFF9",X"FFF7FB",X"F8FFFC",X"FEFFFB",X"FFF9FF",X"FEFFFF",X"E6FEFE",X"5C8EC3",X"0756BF",X"0E74D9",X"0672E1",X"005CC4",X"0A63C7",X"226DD2",X"1B56B4",X"002169",X"000B32",X"27313B",X"070002",X"7F824D",X"DAE062",X"D9D735",X"E5DD56",X"726E27",X"010200",X"000104",X"652A0A",X"ED8F4F",X"F07929",X"FE8A3F",X"F4862F",X"F18314",X"F68B23",X"E28035",X"D38A2B",X"F09745",X"FB8C47",X"FF8339",X"F5781C",X"FC8318",X"FA8416",X"F27D13",X"EE7E01",X"E47C1B",X"E38D52",X"B67E63",X"291715",X"000322",X"073C80",X"2066C8",X"005DD5",X"0C62CF",X"0F61C5",X"146DD5",X"056BD9",X"0666CC",X"2A6FBA",X"2B5689",X"0A0722",X"282A63",X"334390",X"2C509C",X"275EB0",X"185CC1",X"0856C3",X"055BC2",X"126BCF",X"1F5CAD",X"254679",X"0F253C",X"273840",X"0D0014",X"571344",X"9E2C74",X"C01476",X"B5026A",X"C8077A",X"CC0078",X"C60074",X"BA217B",X"6D1B4C",X"1F0415",X"080226",X"16377E",X"1159AE",X"1568C8",X"0052CA",X"0B68E1",X"076DD1",X"0061BF",X"0D6AD4",X"065ECC",X"0458C8",X"0A60CF",X"0862D0",X"0663CB",X"0F6BD2",X"156CD3",X"0F5EC5",X"0B69CD",X"0A62C4",X"2763C3",X"0B3984",X"001743",X"00041B",X"1D1928",X"478383",X"37948C",X"159C8B",X"1AB5A3",X"079F90",X"18AB9B",X"0C9F8D",X"13AC97",X"00907A",X"A4F9F2"),
(X"FFFEFF",X"80DDCB",X"04BD9B",X"2AC9B5",X"0AC9A7",X"00CBA0",X"01BF9B",X"11D2B3",X"1EB999",X"0C4B36",X"000313",X"746B1E",X"ECC319",X"F0D339",X"B4A445",X"000200",X"1B0802",X"1F2521",X"26504E",X"0D5351",X"055657",X"0B6162",X"095E63",X"00545E",X"086260",X"06615C",X"025E59",X"005F5B",X"005D5D",X"0C5C63",X"16555C",X"0A3B42",X"081616",X"000505",X"1F4641",X"58AEA3",X"44D5C8",X"13CDC8",X"0BD7E0",X"07D4E9",X"16DDF2",X"05D0DE",X"00D0D3",X"04D9D5",X"00CEC8",X"0CDAD8",X"0EDEE0",X"03D4D8",X"0EE1EA",X"00D0DB",X"0BDFEA",X"00D5DE",X"00D4D9",X"0FD5D8",X"30D9E0",X"1BABB6",X"00464A",X"00131C",X"000715",X"000109",X"22251E",X"667359",X"889B6E",X"9AB37C",X"82AE5F",X"79AC5D",X"77B464",X"6AAF5F",X"6AB364",X"6CB566",X"76BD6F",X"7EC174",X"6E9674",X"001000",X"000600",X"050500",X"070000",X"3D2D1E",X"715C41",X"917754",X"D39B48",X"E1A44B",X"E79D3C",X"F1952E",X"F88E21",X"FF9A24",X"EB8300",X"F39300",X"DD8837",X"623D10",X"000500",X"820549",X"DB0C76",X"DA1C86",X"C80264",X"EA8ABA",X"FFF8FF",X"FCFDFF",X"FEFCFF",X"FFF9FD",X"FFFCFD",X"F8FFFF",X"F8FFFE",X"FFFBFD",X"F7FFFF",X"C9CACC",X"000103",X"212026",X"152930",X"314560",X"274D7A",X"2C5491",X"3064AF",X"3575BD",X"2C76BF",X"226EBC",X"2161B8",X"2970C8",X"226FC9",X"1A6BC4",X"2273CE",X"1D71D1",X"1770D8",X"106FDB",X"0D6FDC",X"0A6FD7",X"096FD1",X"0A6FCB",X"DADEEA",X"FCFEFF",X"F8FBFF",X"FBFDFC",X"FFFFFD",X"FAFAF8",X"FFFEFF",X"F4F2F5",X"1B1931",X"746718",X"EDD82F",X"E9DD0B",X"F1E90A",X"F0E00E",X"E7D40B",X"ECE308",X"FAE700",X"EFE511",X"DCD32E",X"FFFFB4",X"FFFCF0",X"F7FFF8",X"FBF4FC",X"FFFDFD",X"FEFFFA",X"FEFFFA",X"FEFFFA",X"FEFFFA",X"FEFFFA",X"FEFFFA",X"FEFFFA",X"FEFFFA",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FCFEFB",X"FAFCF9",X"FFFEFF",X"DDC7DC",X"300E02",X"602F33",X"39080E",X"380E12",X"170D0E",X"0C0600",X"050400",X"000107",X"000800",X"001609",X"000700",X"213519",X"1D481A",X"44703D",X"5E8D56",X"53864E",X"A3D8A4",X"8BC18F",X"558E59",X"6DA76D",X"62AC4D",X"5B9549",X"A4C898",X"F5FFEE",X"FDFCFA",X"FEF9FD",X"FFFFFF",X"F3F8F2",X"83AD7F",X"639B52",X"6EA145",X"6FA04E",X"629D5D",X"71A05C",X"84A465",X"668C75",X"47533D",X"13242C",X"00031C",X"9CB0AE",X"F9FEFF",X"FFFBFF",X"FFFFED",X"FCFEFD",X"FDFBFF",X"FFFCFC",X"FFF7FF",X"FBFEFF",X"E3FFF9",X"548EBC",X"0752C9",X"1370CD",X"1A5BC1",X"316AC4",X"2F5C97",X"2F4B61",X"1A272D",X"010000",X"0B0400",X"0B0500",X"A99E2A",X"E3D22A",X"E8DC0C",X"D7D205",X"E8DD1F",X"DFC928",X"4F3F00",X"070A00",X"000200",X"5E3D2E",X"DE9769",X"F6863A",X"FF8124",X"E77C0A",X"F7A02C",X"FA8621",X"FE8325",X"F78008",X"F78407",X"FB8523",X"F47C26",X"EF7812",X"FD8517",X"FA831D",X"EC8D3B",X"E27E28",X"E69858",X"9B7C60",X"30271E",X"0F0704",X"030E20",X"1D4978",X"2A5DB8",X"0A64BA",X"0064C9",X"005DD5",X"076BDB",X"126CCC",X"115BBA",X"0D5DC0",X"124DB1",X"2166B1",X"165CB1",X"2468E3",X"0B5BD8",X"0467C4",X"0866BE",X"175FD5",X"0B68CF",X"0360C8",X"1C66C9",X"2957A4",X"000531",X"00031F",X"4A1948",X"891A66",X"AC1274",X"BA0B74",X"C60778",X"BF006E",X"CA0473",X"C5026B",X"C01973",X"7E0047",X"1F0017",X"0E0018",X"070D31",X"385893",X"3F83D8",X"0164CA",X"0A75DF",X"096CD4",X"0268D4",X"0065CE",X"0063CA",X"0669D1",X"025DC6",X"0B61CE",X"075FCB",X"005DC7",X"146CC5",X"1866B0",X"235C91",X"204162",X"081F31",X"000E14",X"11665F",X"1A9082",X"0DB196",X"08A59A",X"009497",X"14AAA8",X"1CB69E",X"009570",X"10A98D",X"16AA9C",X"0A9292",X"98F5ED"),
(X"FFFCFD",X"7AD7C5",X"0BC4A2",X"25C4B0",X"15D4B2",X"00C89D",X"04C29E",X"07C8A9",X"2DC8A8",X"2E6D58",X"000414",X"685F12",X"EAC117",X"EFD238",X"A19132",X"040905",X"26130D",X"000200",X"1D4745",X"135957",X"095A5B",X"005657",X"03585D",X"075B65",X"005856",X"005A55",X"05615C",X"0A6A66",X"036161",X"04545B",X"16555C",X"1D4E55",X"051313",X"0F2121",X"000C07",X"002B20",X"17A89B",X"2FE9E4",X"07D3DC",X"02CFE4",X"03CADF",X"0CD7E5",X"07DBDE",X"00D3CF",X"02D5CF",X"04D2D0",X"04D4D6",X"09DADE",X"00CFD8",X"0ADDE8",X"06DAE5",X"00D7E0",X"07DEE3",X"09CFD2",X"19C2C9",X"3CCCD7",X"49A8AC",X"3C7F88",X"284553",X"00020A",X"000200",X"000700",X"25380B",X"6E8750",X"89B566",X"7DB061",X"72AF5F",X"73B868",X"69B263",X"63AC5D",X"68AF61",X"7ABD70",X"82AA88",X"658264",X"788571",X"6E6E62",X"170E05",X"0D0000",X"120000",X"190000",X"733B00",X"995C03",X"BE7413",X"EA8E27",X"FF9F32",X"FA8B15",X"FF9E17",X"F69603",X"EA9544",X"6E491C",X"000B02",X"84074B",X"D90A74",X"DA1C86",X"CE086A",X"E888B8",X"FFF8FF",X"FCFDFF",X"FEFCFF",X"FFF9FD",X"FFFDFE",X"F8FFFF",X"F9FFFF",X"FFFBFD",X"F4FFFC",X"C8C9CB",X"0A0B0D",X"141319",X"00050C",X"000722",X"000734",X"00114E",X"00236E",X"003981",X"004089",X"1561AF",X"2363BA",X"1A61B9",X"216EC8",X"2A7BD4",X"2374CF",X"2377D7",X"247DE5",X"207FEB",X"1C7EEB",X"167BE3",X"147ADC",X"1479D5",X"DBDFEB",X"FBFDFF",X"F7FAFF",X"FBFDFC",X"FFFFFD",X"FBFBF9",X"FFFEFF",X"F3F1F4",X"1F1D35",X"6D6011",X"FFEE45",X"FCF01E",X"E7DF00",X"F0E00E",X"FFED24",X"E9E005",X"F4E100",X"F0E612",X"F1E843",X"FDFBB0",X"FFF8EC",X"F7FFF8",X"FFFCFF",X"FFFCFC",X"FEFFFA",X"FEFFFA",X"FEFFFA",X"FEFFFA",X"FEFFFA",X"FEFFFA",X"FEFFFA",X"FEFFFA",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFFFD",X"F3F5F2",X"FFFEFF",X"D5BFD4",X"190000",X"320105",X"48171D",X"451B1F",X"473D3E",X"3B3525",X"0C0B07",X"3C4349",X"4F6455",X"51695C",X"71867F",X"7F9377",X"6F9A6C",X"84B07D",X"7FAE77",X"497C44",X"8CC18D",X"BFF5C3",X"568F5A",X"659F65",X"6FB95A",X"5B9549",X"9DC191",X"F7FFF0",X"FFFFFD",X"F7F2F6",X"FCFCFC",X"F6FBF5",X"88B284",X"619950",X"70A347",X"6D9E4C",X"6DA868",X"78A763",X"4C6C2D",X"052B14",X"020E00",X"0C1D25",X"02162F",X"9DB1AF",X"F8FDFF",X"FFFCFF",X"FFFFEC",X"FEFFFF",X"FEFCFF",X"FFFAFA",X"FFF8FF",X"F4F7FF",X"E4FFFA",X"5892C0",X"0B56CD",X"1673D0",X"1D5EC4",X"124BA5",X"001A55",X"000B21",X"00050B",X"010000",X"8D8669",X"BFB97B",X"DFD460",X"DDCC24",X"DDD101",X"DDD80B",X"D4C90B",X"F7E140",X"BFAF57",X"000200",X"000604",X"190000",X"A96234",X"F08034",X"FF781B",X"E97E0C",X"E08915",X"FB8722",X"FD8224",X"F78008",X"F98609",X"F7811F",X"FB832D",X"F67F19",X"EA7204",X"EA730D",X"F99A48",X"EC8832",X"AC5E1E",X"3E1F03",X"170E05",X"090100",X"000113",X"022E5D",X"1F52AD",X"126CC2",X"1177DC",X"005BD3",X"005ECE",X"0D67C7",X"1B65C4",X"0050B3",X"0A45A9",X"1156A1",X"1056AB",X"1559D4",X"1464E1",X"0C6FCC",X"0058B0",X"1D65DB",X"126FD6",X"0764CC",X"1660C3",X"2B59A6",X"22416D",X"000723",X"1D001B",X"640041",X"A70D6F",X"C1127B",X"BD006F",X"C60675",X"CA0473",X"CD0A73",X"B30C66",X"BE3B87",X"401438",X"1E0928",X"00062A",X"001B56",X"1A5EB3",X"0C6FD5",X"0068D2",X"1275DD",X"005CC8",X"0068D1",X"0066CD",X"0061C9",X"045FC8",X"055BC8",X"025AC6",X"0865CF",X"1E76CF",X"1967B1",X"00356A",X"00092A",X"152C3E",X"154046",X"429790",X"259B8D",X"009C81",X"10ADA2",X"0DA5A8",X"049A98",X"17B199",X"10AC87",X"11AA8E",X"10A496",X"008585",X"92EFE7"),
(X"FEFCFD",X"79DAC6",X"00BF97",X"1BC7AD",X"0AC9A7",X"09C7A1",X"06BE9C",X"05C7A5",X"2BD3B9",X"288884",X"00050C",X"3E2F1A",X"E0B950",X"D1BD4A",X"261C03",X"100000",X"400F00",X"2A0700",X"070000",X"1C3637",X"1E5657",X"0E5A58",X"106260",X"0B5C5D",X"055B6A",X"025962",X"025C5C",X"086761",X"02625E",X"005B5A",X"055E62",X"0B5E64",X"0D5B5D",X"002024",X"001420",X"050012",X"030015",X"517C8C",X"55D1CF",X"25E0CF",X"0BD1DA",X"00CCD7",X"07D7E4",X"01D3E4",X"02D1E1",X"00CAD7",X"07D8DC",X"05DAD8",X"00D4D6",X"0BDCE1",X"0AD2DF",X"0DD6E6",X"00CFDC",X"05D9E5",X"00D3DC",X"0AD6DF",X"0CD4E3",X"20D4E3",X"2DC3D4",X"0E8492",X"001F29",X"001519",X"071516",X"060000",X"3C442C",X"728361",X"82A374",X"8CBA7C",X"80B56F",X"7AAF67",X"79AB64",X"74A15E",X"6AB269",X"79BB73",X"7EBA74",X"7AB072",X"497947",X"3B613A",X"213C1B",X"000800",X"000204",X"0B0A05",X"0A0000",X"3D2E0D",X"786837",X"9B7E42",X"D29D57",X"DF974D",X"E6A97C",X"7D4536",X"0A0000",X"811048",X"D41879",X"DF1585",X"D80067",X"EB89B0",X"FFF6FF",X"FCFDFF",X"FEFEFF",X"FFFBFE",X"FFFDFE",X"F9FFFF",X"FBFFFF",X"FFFAFD",X"FFF6FF",X"C3E1E1",X"006A4F",X"005D55",X"003A36",X"001B24",X"000A13",X"000F19",X"040003",X"0C0109",X"040005",X"000B0A",X"13000F",X"00050F",X"00040B",X"001015",X"001549",X"052057",X"0F2D69",X"153977",X"18407E",X"1B4380",X"204780",X"234B7F",X"E2E4F0",X"FBFEFF",X"F6FAFD",X"FBFDFC",X"FFFFFD",X"FCFCFA",X"FFFEFF",X"F2F0F3",X"252736",X"504C1F",X"C2BA69",X"CDCA69",X"DFDC69",X"E2D660",X"E5DC67",X"DFE962",X"EFE75E",X"E4E065",X"F2E77E",X"FDFFD0",X"FFFEF8",X"F0FFF4",X"FBFFFF",X"F4FDF8",X"FEFEFC",X"FEFEFC",X"FEFEFC",X"FEFEFC",X"FEFEFC",X"FEFEFC",X"FEFEFC",X"FEFEFC",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEF7FE",X"FFFEFF",X"EFF4EE",X"CEDADA",X"0A2700",X"4C7040",X"74A16A",X"7CAE73",X"7FA56C",X"6C9350",X"5B8546",X"7EAF78",X"6EA967",X"69A75E",X"76AE6D",X"6EA065",X"618955",X"588149",X"5E8A4F",X"517D42",X"527F48",X"A9D8A2",X"8ABB83",X"57894C",X"5F8B50",X"527346",X"97A98F",X"F5FBF1",X"FFFEFF",X"FEFCFD",X"FEFFFD",X"F8FFF8",X"7BA07F",X"6AA064",X"719F70",X"699266",X"7EA996",X"5B6F70",X"000100",X"000028",X"00104D",X"1B3F97",X"13369E",X"94B0E2",X"F5FDFF",X"FFFDFF",X"FDF9F8",X"FCFCFF",X"FEFFFD",X"FBFBF3",X"FFFDFF",X"FEFFFF",X"EAFDFF",X"6383C0",X"2852B8",X"215B9B",X"1E3352",X"001119",X"0C1206",X"0F0800",X"231400",X"9B8C0B",X"E3D625",X"EADE18",X"DCCC00",X"F2CE06",X"F3CB11",X"DCC60E",X"DBD40A",X"DFD60B",X"DED230",X"8A8414",X"41371E",X"483A37",X"0B0001",X"986959",X"E88B50",X"F18D2B",X"EC831A",X"FF7828",X"FF7D13",X"FD7D00",X"F88200",X"F58508",X"E97909",X"FF9333",X"E3813A",X"DB8A5F",X"A27A56",X"5A3B38",X"130000",X"150000",X"483D00",X"838732",X"141A00",X"01000E",X"141E5B",X"1659A8",X"0A63C9",X"0A58C4",X"2B7AD7",X"1C5AA7",X"3B4D7B",X"7D717B",X"7E6E7B",X"7B616C",X"5E5769",X"1D4076",X"1758BE",X"155EE1",X"045AD3",X"0065C9",X"0C74E5",X"026EDB",X"0062D2",X"0C5FD7",X"2470DE",X"00357D",X"00051C",X"160300",X"41043F",X"8A226D",X"C21E7F",X"D10576",X"CF006F",X"CE0F79",X"BF0F72",X"C31979",X"B01678",X"670C51",X"320D2F",X"10000E",X"030015",X"40688C",X"438BD3",X"004CB4",X"104FB6",X"0D5AC6",X"005ACC",X"0B6BE3",X"0461D8",X"1062D0",X"0C54B6",X"195CB5",X"1E5385",X"0B2A59",X"000128",X"000B1E",X"00534E",X"22AF9C",X"1BBDA8",X"09AB9C",X"109A8A",X"12A68C",X"0EAE8A",X"0CB58C",X"05AF88",X"16BA98",X"059F85",X"0EA08B",X"1C8769",X"B2F6DD"),
(X"FDFBFC",X"7ADBC7",X"00BB93",X"1BC7AD",X"02C19F",X"0AC8A2",X"04BC9A",X"02C4A2",X"21C9AF",X"389894",X"02161D",X"0D0000",X"D9B249",X"C4B03D",X"0C0200",X"251305",X"A37252",X"8B6854",X"080000",X"001011",X"003637",X"095553",X"015351",X"095A5B",X"055B6A",X"065D66",X"005A5A",X"005E58",X"005F5B",X"005F5E",X"065F63",X"03565C",X"0F5D5F",X"256064",X"0F2733",X"050012",X"0C071E",X"000B1B",X"169290",X"17D2C1",X"14DAE3",X"06D2DD",X"0ADAE7",X"06D8E9",X"02D1E1",X"02D0DD",X"06D7DB",X"00CBC9",X"09E0E2",X"01D2D7",X"07CFDC",X"12DBEB",X"00C9D6",X"0ADEEA",X"0CDFE8",X"00CAD3",X"11D9E8",X"16CAD9",X"2CC2D3",X"45BBC9",X"469AA4",X"002B2F",X"000405",X"100708",X"000500",X"000B00",X"416233",X"719F61",X"7AAF69",X"84B971",X"77A962",X"77A461",X"6BB36A",X"6DAF67",X"68A45E",X"70A668",X"89B987",X"8DB38C",X"839E7D",X"617154",X"2D3537",X"2E2D28",X"1D1200",X"140500",X"150500",X"210400",X"582300",X"B56D23",X"A36639",X"622A1B",X"0A0000",X"800F47",X"D71B7C",X"DF1585",X"D50064",X"EC8AB1",X"FFF6FF",X"FBFCFF",X"FEFEFF",X"FFFBFE",X"FFFDFE",X"F9FFFF",X"FBFFFF",X"FFFBFE",X"FFF0F9",X"CAE8E8",X"14A085",X"44A8A0",X"3F9894",X"47737C",X"2D525B",X"2A4C56",X"0B060A",X"070004",X"050006",X"000807",X"574253",X"A8AFB9",X"9DACB3",X"9FB4B9",X"90A7DB",X"92ADE4",X"93B1ED",X"90B4F2",X"8BB3F1",X"8AB2EF",X"8DB4ED",X"90B8EC",X"EBEDF9",X"FCFFFF",X"F7FBFE",X"FBFDFC",X"FEFEFC",X"FDFDFB",X"FFFEFF",X"F2F0F3",X"3A3C4B",X"080400",X"140C00",X"2E2B00",X"6D6A00",X"685C00",X"5C5300",X"89930C",X"9D950C",X"848005",X"8E831A",X"EBEDBE",X"FFFDF7",X"EFFFF3",X"FBFFFF",X"F9FFFD",X"FEFEFC",X"FEFEFC",X"FEFEFC",X"FEFEFC",X"FEFEFC",X"FEFEFC",X"FEFEFC",X"FEFEFC",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FFFCFF",X"FEFCFD",X"FCFFFB",X"C6D2D2",X"7B9862",X"80A474",X"90BD86",X"6A9C61",X"7AA067",X"729956",X"7EA869",X"78A972",X"619C5A",X"68A65D",X"5F9756",X"90C287",X"B2DAA6",X"B4DDA5",X"AEDA9F",X"B5E1A6",X"A8D59E",X"B9E8B2",X"C7F8C0",X"9ED093",X"B0DCA1",X"A9CA9D",X"CCDEC4",X"F9FFF5",X"FEFCFD",X"FCFAFB",X"FBFDFA",X"EDF4ED",X"98BD9C",X"70A66A",X"7BA97A",X"4E774B",X"001300",X"021617",X"000100",X"16153F",X"2F4F8C",X"4064BC",X"2346AE",X"93AFE1",X"F8FFFF",X"FFFDFF",X"FBF7F6",X"FBFBFF",X"FEFFFD",X"FDFDF5",X"FFFDFF",X"FEFFFF",X"EBFEFF",X"6686C3",X"123CA2",X"0E4888",X"000322",X"000810",X"000500",X"60593C",X"D2C37E",X"D9CA49",X"D7CA19",X"D0C400",X"ECDC0D",X"F3CF07",X"EFC70D",X"DDC70F",X"E9E218",X"D2C900",X"DCD02E",X"DBD565",X"9C9279",X"2C1E1B",X"0E0004",X"3E0F00",X"CB6E33",X"E37F1D",X"F28920",X"FE7121",X"FF841A",X"F37300",X"FA8400",X"F18104",X"F88818",X"FF9232",X"DD7B34",X"A35227",X"290100",X"160000",X"110000",X"755E35",X"C0B55C",X"D0D47F",X"717755",X"02000F",X"06104D",X"003584",X"0760C6",X"1664D0",X"0352AF",X"2765B2",X"7E90BE",X"9E929C",X"A393A0",X"B49AA5",X"948D9F",X"6386BC",X"2162C8",X"145DE0",X"146AE3",X"016BCF",X"0169DA",X"026EDB",X"0367D7",X"0A5DD5",X"1561CF",X"1E5EA6",X"19334A",X"140100",X"260024",X"640047",X"AF0B6C",X"D20677",X"D50275",X"BD0068",X"BC0C6F",X"B60C6C",X"A60C6E",X"680D52",X"532E50",X"1D081B",X"020014",X"083054",X"266EB6",X"1663CB",X"1A59C0",X"0956C2",X"0762D4",X"0767DF",X"004FC6",X"0658C6",X"1E66C8",X"1E61BA",X"003466",X"000433",X"15244B",X"32586B",X"338E89",X"25B29F",X"0FB19C",X"02A495",X"0E9888",X"009278",X"03A37F",X"0CB58C",X"00A881",X"0BAF8D",X"0CA68C",X"1EB09B",X"0E795B",X"B3F7DE"),
(X"FCFAFB",X"7AD1BE",X"03C69A",X"13CBA9",X"0ECDAB",X"0DC0A0",X"0FBEA1",X"00BE9D",X"11CDB4",X"2AB8AA",X"0D4A42",X"110012",X"A6986B",X"776130",X"0A0C18",X"5C2500",X"F28A29",X"CD7A34",X"270000",X"140000",X"0A000D",X"16272F",X"2C6157",X"0B5B42",X"025156",X"0A5B5F",X"06595F",X"055D61",X"045F60",X"005F5D",X"006258",X"005D51",X"115F6C",X"00585C",X"0B615E",X"08403F",X"00040B",X"111520",X"00070C",X"255957",X"43B7AE",X"3CC5BD",X"1FC5C1",X"12CFD3",X"12D8E5",X"0FD2E6",X"04C2DA",X"0EC8E1",X"07D8D3",X"06D2D1",X"05CFD3",X"0DD8DF",X"08DBE2",X"01D8DD",X"00D7DC",X"0CE1E5",X"08D2E0",X"0FD7E4",X"03C8D0",X"13D3D6",X"19C7C6",X"2EC0BD",X"0E817E",X"002B2B",X"00090D",X"03161C",X"000209",X"000102",X"4F5748",X"708660",X"7FA76B",X"83B76D",X"81AA64",X"78AA61",X"73B168",X"62AD68",X"65B673",X"61A967",X"76AD69",X"8DB76F",X"87B97A",X"7BB674",X"6AA66A",X"133E11",X"001300",X"000400",X"000202",X"000705",X"000700",X"200806",X"0C0003",X"800E42",X"D71377",X"EF138E",X"D90065",X"EB85AA",X"FFF4FE",X"FCFBFF",X"FDFEFF",X"FFFCFE",X"FFFCFE",X"FBFFFF",X"FCFFFF",X"FFFBFE",X"F8FFFF",X"B1F5E8",X"02AB8A",X"1CB8A3",X"27BAA8",X"0BC59C",X"22B38A",X"29BB8A",X"09987C",X"188C79",X"188474",X"007454",X"6B9999",X"E7FFFF",X"F9FDFF",X"FDFAFF",X"FFFDFF",X"FFFDFF",X"FEFFFF",X"FBFFFF",X"F9FFFF",X"FBFFFF",X"FBFFFF",X"FCFFFF",X"F6F9FE",X"FCFFFF",X"FBFDFC",X"FCFEFB",X"FDFDFB",X"FDFDFB",X"FFFEFF",X"F3F1F4",X"233040",X"070B0A",X"120F18",X"010010",X"080000",X"170100",X"0A0000",X"040D00",X"02020E",X"000004",X"170500",X"E2E1E6",X"FFFAFF",X"FBFFF6",X"FFF9F9",X"FEFAF1",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"F7F6FC",X"FEFCFD",X"FCFFF8",X"C6DED0",X"5F974C",X"5DA156",X"60A555",X"7DBC6B",X"6BA25E",X"75AD64",X"679F54",X"65A15B",X"6FAE67",X"66A650",X"649A4F",X"C7F0CE",X"FEFDFF",X"FFFFFF",X"FCFCFA",X"F3F5F4",X"FEFFFF",X"FCFDFF",X"F3F4F6",X"FCFFFD",X"F9FFF6",X"F9FFF5",X"FEFFFA",X"FEFCFD",X"FBF6FA",X"FFFEFF",X"FEFFFD",X"FAFFF9",X"AEAE96",X"394A28",X"3F4150",X"000010",X"00002E",X"00014A",X"0F4470",X"1E65BF",X"1F67D3",X"1B67D5",X"0247C0",X"7EADE5",X"F1FFFA",X"FFFFF1",X"FFFFF3",X"F8FDFF",X"FBFEFF",X"FCFBFF",X"FFFDFF",X"F2F2EA",X"FCFFFF",X"878BB1",X"000015",X"22301F",X"040100",X"0F1000",X"7F8100",X"DBD833",X"E2DC24",X"D6CE07",X"D9D10A",X"D9D011",X"D0C500",X"E5D900",X"E0D700",X"DACF13",X"E3CF16",X"E5C80A",X"F4DB4D",X"C6B871",X"49432B",X"1A0000",X"310617",X"220000",X"2E0000",X"A5764C",X"DA9753",X"F68340",X"ED821A",X"EB7714",X"EB7D1C",X"E78D2D",X"DF8D43",X"B26841",X"593424",X"000300",X"140000",X"130800",X"C1BC44",X"D3D045",X"E1DB69",X"959058",X"39393B",X"000026",X"001363",X"0E4EA6",X"1B68D4",X"1269DC",X"1258AE",X"7E7796",X"DB7F5A",X"F1781B",X"E77419",X"ED7224",X"F77D34",X"DF7F43",X"9F7370",X"354C92",X"0F62C2",X"006DC0",X"0A5EE2",X"0564CE",X"036BC2",X"0060BC",X"005FC8",X"1C7CE2",X"2463B2",X"00164E",X"110D2E",X"27103A",X"661758",X"AB116F",X"CA0674",X"C90573",X"C60673",X"F32E9A",X"D92265",X"BD0964",X"AB1E7A",X"581349",X"13000C",X"050110",X"000738",X"2861B0",X"1761CC",X"0050BA",X"0E67CF",X"0A61C2",X"1D65B9",X"265D9E",X"406997",X"2A4B6C",X"000B15",X"003A39",X"007364",X"1AA892",X"14A892",X"0CA18E",X"1FBCAB",X"00A694",X"009E7C",X"11AA8C",X"1CAC95",X"089B89",X"10A899",X"17A494",X"34A393",X"419888",X"0C3120",X"D2D3CD"),
(X"FFFEFF",X"7CD3C0",X"00C397",X"17CFAD",X"0BCAA8",X"10C3A3",X"11C0A3",X"04C3A2",X"0DC9B0",X"1AA89A",X"00352D",X"0E000F",X"67592C",X"513B0A",X"00000B",X"7D461F",X"EC8423",X"D6833D",X"915F3C",X"170000",X"140917",X"000D15",X"02372D",X"0C5C43",X"0D5C61",X"0D5E62",X"04575D",X"055D61",X"076263",X"005F5D",X"006359",X"016559",X"0B5966",X"035C60",X"0C625F",X"28605F",X"23343B",X"010510",X"031C21",X"00100E",X"00433A",X"129B93",X"2FD5D1",X"20DDE1",X"03C9D6",X"0BCEE2",X"0FCDE5",X"19D3EC",X"00CEC9",X"09D5D4",X"08D2D6",X"01CCD3",X"0BDEE5",X"00D5DA",X"00D3D8",X"0BE0E4",X"0FD9E7",X"0CD4E1",X"11D6DE",X"11D1D4",X"23D1D0",X"2CBEBB",X"48BBB8",X"419B9B",X"30494D",X"00080E",X"000209",X"0A0E0F",X"010900",X"000B00",X"4C7438",X"6A9E54",X"89B26C",X"82B46B",X"79B76E",X"64AF6A",X"5DAE6B",X"71B977",X"72A965",X"739D55",X"80B273",X"71AC6A",X"86C286",X"85B083",X"728571",X"5F645E",X"424848",X"15211F",X"000700",X"130000",X"0D0004",X"841246",X"D81478",X"F0148F",X"D50061",X"E882A7",X"FEF2FC",X"FBFAFF",X"FDFEFF",X"FFFCFE",X"FFFCFE",X"FAFFFE",X"FBFFFE",X"FFFBFE",X"F4FFFB",X"ABEFE2",X"01AA89",X"1DB9A4",X"24B7A5",X"04BE95",X"1EAF86",X"21B382",X"22B195",X"3EB29F",X"3CA898",X"0FA484",X"81AFAF",X"DCFEFF",X"F9FDFF",X"FFFDFF",X"FFFDFF",X"FFFCFF",X"FBFCFF",X"F7FCFF",X"F5FCFF",X"F7FBFF",X"F6FAFF",X"F6F9FF",X"FCFFFF",X"FCFFFF",X"FDFFFE",X"FDFFFC",X"FCFCFA",X"FEFEFC",X"FFFEFF",X"F4F2F5",X"323F4F",X"000100",X"0B0811",X"0D081C",X"0F0402",X"200A00",X"160900",X"0E1706",X"191925",X"18171C",X"0E0000",X"EAE9EE",X"FFF7FF",X"F7FFF2",X"FFFBFB",X"FFFFF6",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FAF8F9",X"FBFFF7",X"CBE3D5",X"5D954A",X"6EB267",X"5EA353",X"6FAE5D",X"679E5A",X"679F56",X"659D52",X"68A45E",X"67A65F",X"65A54F",X"6AA055",X"BEE7C5",X"FFFEFF",X"FAFAFC",X"FFFFFD",X"FAFCFB",X"FAFBFF",X"FEFFFF",X"F9FAFC",X"FCFFFD",X"F5FFF2",X"FBFFF7",X"FFFFFB",X"FFFDFE",X"FDF8FC",X"FDFBFC",X"FAFCF9",X"F3F8F2",X"97977F",X"011200",X"030514",X"030214",X"253765",X"3757A0",X"2F6490",X"135AB4",X"175FCB",X"1460CE",X"074CC5",X"79A8E0",X"EAFEF3",X"FFFEEF",X"FFFFF4",X"F7FCFF",X"FCFFFF",X"FAF9FF",X"F6F1F5",X"FFFFF8",X"F4F7FF",X"61658B",X"000015",X"000800",X"2A2718",X"A4A55F",X"D9DB56",X"D7D42F",X"C8C20A",X"D8D009",X"CCC400",X"E2D91A",X"E8DD11",X"DBCF00",X"E3DA01",X"D9CE12",X"DDC910",X"FBDE20",X"C6AD1F",X"372900",X"090300",X"3B1D1B",X"3D1223",X"410E1F",X"45100A",X"260000",X"C4813D",X"FB8845",X"E67B13",X"FD8926",X"F88A29",X"CB7111",X"9F4D03",X"4E0400",X"1F0000",X"030900",X"988354",X"C3B869",X"C9C44C",X"D3D045",X"AAA432",X"110C00",X"030305",X"090B31",X"2750A0",X"2767BF",X"1360CC",X"0960D3",X"0E54AA",X"87809F",X"DA7E59",X"FF8629",X"EF7C21",X"EB7022",X"F67C33",X"D37337",X"BF9390",X"556CB2",X"095CBC",X"0071C4",X"0053D7",X"0B6AD4",X"1A82D9",X"056ECA",X"0066CF",X"0868CE",X"2F6EBD",X"39568E",X"2E2A4B",X"37204A",X"8E3F80",X"AC1270",X"BF0069",X"C70371",X"B70064",X"D20D79",X"C30C4F",X"BF0B66",X"AE217D",X"712C62",X"190212",X"0C0817",X"000536",X"003685",X"226CD7",X"0A5DC7",X"035CC4",X"136ACB",X"145CB0",X"003071",X"00103E",X"001132",X"365E68",X"539B9A",X"2DA091",X"23B19B",X"0CA08A",X"0BA08D",X"0EAB9A",X"04AB99",X"03A785",X"08A183",X"12A28B",X"1FB2A0",X"029A8B",X"129F8F",X"239282",X"005343",X"000F00",X"CECFC9"),
(X"FFFEFF",X"90CABC",X"09AE86",X"1DCDA9",X"00C29C",X"0FC6A7",X"0EBDA0",X"0AC3A3",X"00C0A2",X"18D9A2",X"128371",X"00060B",X"080000",X"120807",X"120000",X"C86E20",X"F37A05",X"FF851D",X"F27E27",X"B85D17",X"2B0000",X"150100",X"0C0C04",X"1B1F2A",X"1B4F4D",X"1C5858",X"0F5555",X"075756",X"0A5C58",X"065B54",X"0A6057",X"0E645B",X"0E5D62",X"015D5A",X"006357",X"006454",X"086457",X"064441",X"02232A",X"011120",X"0F0007",X"040B11",X"20514D",X"4DAA9F",X"49CFC4",X"25CCC5",X"07C7C8",X"00CFD5",X"00D0D4",X"05D6DD",X"09D5DE",X"00CAD5",X"05D1DC",X"05D4DC",X"04D5DA",X"00CED3",X"01D2D7",X"0BDEE5",X"04D8E3",X"04DDE6",X"00D6DF",X"02D8E0",X"04D5DC",X"0AD5DC",X"13C8CF",X"0FACB1",X"057B7B",X"001615",X"000D09",X"011513",X"000304",X"020A0D",X"4E5F55",X"6D8168",X"94B280",X"8FBA75",X"70A65A",X"71AE61",X"78B46A",X"72AB64",X"62B25D",X"62AA54",X"68A651",X"80B968",X"75AF63",X"87C37D",X"81BA73",X"70A85F",X"4A6D4D",X"121814",X"00000B",X"861B53",X"D8157B",X"E8178E",X"C60064",X"EE7CB0",X"FFEFFB",X"FCF9FF",X"FBFFFF",X"FFFDFE",X"FFFBFD",X"FBFFFE",X"FDFFFE",X"FFFAFD",X"FFFEFF",X"C5E9DF",X"04A579",X"27B197",X"00C29B",X"00BC96",X"00BB96",X"0AB593",X"00B995",X"0DAD91",X"0DA68A",X"02AC88",X"6CC4B6",X"E4FEFD",X"FFF6FF",X"FFF1F6",X"FFFDF8",X"FFFDF6",X"FFFFF5",X"FFFFF6",X"FFFFF6",X"FFFFF8",X"FFFFFB",X"FFFFFD",X"FEFFFF",X"FEFFFF",X"FEFFFD",X"FFFFFD",X"FDFDFB",X"FEFEFE",X"FFFEFF",X"F4F2F5",X"3F3734",X"1E0000",X"500315",X"4E0016",X"560006",X"500000",X"490004",X"490014",X"240000",X"2D0004",X"2A0000",X"EDE2DE",X"FFFDFF",X"FFFFF4",X"FFFCFF",X"FFFBFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"F9FEFF",X"F9F9F7",X"FFFFF4",X"CCE1D0",X"588C41",X"73B168",X"71A35C",X"789B57",X"70B65E",X"60A353",X"71B457",X"6AAC54",X"599A48",X"69AA46",X"6FA34E",X"BBDDC4",X"F5F5FF",X"FEFFFF",X"FEFFFF",X"FCFDFF",X"FDFDFF",X"FFFDFF",X"FDFCFF",X"FDFCFF",X"FFFBFF",X"FFFDFF",X"FFFDFF",X"FFFDFF",X"FFFEFF",X"FEFCFD",X"FDFBFC",X"FFFEFF",X"A5AABD",X"00072E",X"053780",X"1A529F",X"2371D3",X"0D64D7",X"0A66CB",X"0D71ED",X"0368EA",X"0A74DA",X"065EC8",X"6CA8DC",X"E7FBF9",X"FFF9FD",X"FFFEFD",X"F5FFF4",X"FAFDF4",X"FCFEF1",X"FFFFF6",X"F4F1E8",X"FFFBFF",X"7B7269",X"100700",X"6D5D0F",X"C5BD1C",X"DCD127",X"DED113",X"DDCB05",X"E5CF19",X"E0C820",X"EDDA1C",X"E0D400",X"E7D00E",X"E4D210",X"DFD418",X"CAC418",X"DED450",X"B6A555",X"483B19",X"070300",X"340000",X"660000",X"C62324",X"B21121",X"62000F",X"572232",X"412318",X"B98E6B",X"F2B073",X"CA854C",X"96624A",X"1C0814",X"040000",X"0E0300",X"6A6700",X"95A61A",X"E3CF30",X"ECDD42",X"DFD750",X"C5BF67",X"282A12",X"000223",X"002869",X"18539F",X"0F6EDC",X"1267D2",X"196ADF",X"0464DD",X"044DA9",X"A086A1",X"F88250",X"FD740A",X"E17B0F",X"FE8C2C",X"FF7A1B",X"FF802D",X"CF7B63",X"7776B0",X"074CB4",X"0A6FDB",X"1966CE",X"1664D0",X"0E5ECD",X"0F61CD",X"2477D7",X"266AB5",X"284D84",X"343C6A",X"1E002D",X"25002F",X"7B286E",X"A51672",X"C40974",X"C5016D",X"BF0269",X"C00A6E",X"B90D85",X"AA2171",X"702442",X"1E0815",X"04082D",X"000045",X"032C86",X"0F54B1",X"0865CF",X"166BC6",X"1C5FA6",X"2B598A",X"0E2946",X"00091B",X"000E18",X"2D444A",X"3CA793",X"2AA48F",X"1DA893",X"0CA48F",X"15B19C",X"008F7A",X"00987E",X"1AB798",X"00A782",X"17B9A2",X"00958C",X"29AEA9",X"44B2A9",X"307B76",X"10323C",X"303650",X"000727",X"CBD0E6"),
(X"FFFEFF",X"83BDAF",X"09AE86",X"15C5A1",X"06CAA4",X"06BD9E",X"0CBB9E",X"00B999",X"00C1A3",X"0DCE97",X"3BAC9A",X"001419",X"190F05",X"070000",X"47311A",X"D17729",X"F87F0A",X"F2770F",X"EE7A23",X"DB803A",X"A5703A",X"54401F",X"010100",X"00030E",X"002927",X"145050",X"185E5E",X"0A5A59",X"035551",X"00554E",X"085E55",X"0B6158",X"07565B",X"015D5A",X"00675B",X"006A5A",X"046053",X"215F5C",X"294A51",X"263645",X"1C0814",X"01080E",X"00130F",X"003C31",X"0F958A",X"1BC2BB",X"10D0D1",X"05D4DA",X"00D3D7",X"05D6DD",X"08D4DD",X"08D4DF",X"08D4DF",X"02D1D9",X"00CFD4",X"04D5DA",X"02D3D8",X"00CDD4",X"01D5E0",X"03DCE5",X"03DCE5",X"03D9E1",X"09DAE1",X"07D2D9",X"18CDD4",X"2BC8CD",X"47BDBD",X"5AA4A3",X"38615D",X"001311",X"00090A",X"000205",X"000900",X"000900",X"365422",X"719C57",X"85BB6F",X"73B063",X"81BD73",X"71AA63",X"62B25D",X"6FB761",X"77B560",X"6EA756",X"72AC60",X"70AC66",X"6DA65F",X"87BF76",X"8CAF8F",X"232925",X"01030F",X"891E56",X"D00D73",X"EA1990",X"CC016A",X"ED7BAF",X"FFEFFB",X"FBF8FF",X"FBFFFF",X"FFFDFE",X"FFFBFD",X"FAFEFD",X"FDFFFE",X"FFFAFD",X"FFFDFE",X"C1E5DB",X"009C70",X"26B096",X"00C59E",X"00C39D",X"03C5A0",X"10BB99",X"00B894",X"0BAB8F",X"1DB69A",X"00A884",X"5BB3A5",X"E3FDFC",X"FFF4FD",X"FFF8FD",X"FFFEF9",X"FFFEF7",X"FFFFF6",X"FFFFF6",X"FFFFF6",X"FFFFF8",X"FFFFFB",X"FFFEFC",X"FEFFFF",X"FCFEFD",X"FEFFFD",X"FFFFFD",X"FEFEFC",X"FFFFFF",X"FFFEFF",X"F4F2F5",X"413936",X"2D0500",X"7B2E40",X"781D40",X"872937",X"7B1721",X"7C1C37",X"6C1937",X"501B2B",X"4E1F25",X"460C00",X"E9DEDA",X"FFFDFF",X"FBFDF0",X"FFFCFF",X"FFFAFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FBFFFF",X"FDFDFB",X"FEFFF3",X"CDE2D1",X"5D9146",X"6BA960",X"6B9D56",X"7C9F5B",X"62A850",X"64A757",X"5FA245",X"69AB53",X"74B563",X"6BAC48",X"689C47",X"C8EAD1",X"FEFEFF",X"F7F8FD",X"FEFFFF",X"FDFEFF",X"FEFEFF",X"FEFCFF",X"FFFEFF",X"FEFDFF",X"FFFBFF",X"FFFDFF",X"FFFCFF",X"FEFCFF",X"FFFEFF",X"FEFCFD",X"FBF9FA",X"FFFEFF",X"CBD0E3",X"0A3158",X"4375BE",X"2961AE",X"1563C5",X"075ED1",X"0662C7",X"0367E3",X"0267E9",X"0A74DA",X"025AC4",X"68A4D8",X"EFFFFF",X"FFFDFF",X"FFFEFD",X"F7FFF6",X"FDFFF7",X"FCFEF1",X"FFFEF5",X"FFFEF5",X"FDF5FF",X"746B62",X"807732",X"D8C87A",X"DED635",X"DACF25",X"D0C305",X"E6D40E",X"DBC50F",X"E1C921",X"E3D012",X"E0D400",X"E2CB09",X"E4D210",X"DED317",X"DAD428",X"B6AC28",X"3D2C00",X"0E0100",X"130F06",X"460A0A",X"92201F",X"BD1A1B",X"B41323",X"8F213C",X"400B1B",X"160000",X"5A2F0C",X"C28043",X"7B3600",X"2B0000",X"13000B",X"040000",X"9F945C",X"D2CF5C",X"CBDC50",X"D4C021",X"DFD035",X"B6AE27",X"352F00",X"010300",X"15294A",X"265293",X"2E69B5",X"106FDD",X"0459C4",X"1F70E5",X"0A6AE3",X"014AA6",X"9A809B",X"F7814F",X"F76E04",X"EC861A",X"EF7D1D",X"F36E0F",X"F26E1B",X"D27E66",X"5A5993",X"1A5FC7",X"0B70DC",X"0C59C1",X"1563CF",X"0656C5",X"1668D4",X"1568C8",X"0E529D",X"00144B",X"00002D",X"1F002E",X"52275C",X"620F55",X"A1126E",X"C40974",X"CA0672",X"C2056C",X"C81276",X"B60A82",X"9B1262",X"450017",X"0F0006",X"04082D",X"374890",X"315AB4",X"2E73D0",X"005AC4",X"1065C0",X"2669B0",X"002455",X"000825",X"000618",X"2B3D47",X"374E54",X"0D7864",X"28A28D",X"1EA994",X"11A994",X"019D88",X"009782",X"12AC92",X"07A485",X"06B08B",X"00A28B",X"0BA198",X"1CA19C",X"319F96",X"002F2A",X"000B15",X"252B45",X"000F2F",X"D1D6EC"),
(X"FFFDFE",X"879A98",X"229578",X"27C5A4",X"00C69F",X"09CBA9",X"09BDA0",X"09BC9E",X"03BEA3",X"02D69B",X"33C3AA",X"1D614A",X"100005",X"010002",X"B06522",X"E9780E",X"FF6E00",X"F67100",X"FA8408",X"F4810C",X"F78522",X"DB762E",X"621B00",X"300400",X"0F0705",X"0D1B1B",X"295351",X"145750",X"0A574D",X"085952",X"0A5B5E",X"055762",X"005554",X"0B5A5E",X"0B5057",X"0F595C",X"0C6261",X"025E5B",X"0A605F",X"0D5B5D",X"085251",X"002223",X"001215",X"000107",X"00060C",X"1C403E",X"409085",X"4CBBAA",X"32C3D6",X"25C7D6",X"12CED9",X"06D5DD",X"01D5E0",X"00CBDA",X"09C7DD",X"1ACFEA",X"00CFD1",X"00D5DA",X"00D0DB",X"02D4E3",X"02D1E1",X"09D8E8",X"04D6E5",X"09DDE9",X"00D0CA",X"04D4D4",X"0FD8DF",X"18D2DF",X"1DC5D2",X"1BABB6",X"007B82",X"004C4E",X"000E09",X"001310",X"000100",X"060000",X"535047",X"6A7A60",X"7EA377",X"83B67B",X"82AA6E",X"7CA664",X"7DB065",X"75B262",X"79BA68",X"79B464",X"77A658",X"91B366",X"79A66D",X"2E3428",X"090013",X"821453",X"DC1477",X"EF1F8F",X"B50064",X"E177B9",X"FFEAF9",X"FFFBFF",X"F8FEFE",X"FFFEFF",X"FFFBFD",X"FEFFFF",X"FCFEFD",X"FFFCFE",X"FFF9FF",X"DCE7E3",X"366F5E",X"32A98D",X"1BBB9F",X"00C1A2",X"09BBA3",X"0FB59F",X"04C5A6",X"0CBDA3",X"11BFA4",X"13AB94",X"38C1A7",X"DDFFFF",X"FFFDFF",X"F4FDF8",X"FFFAFF",X"FFFCFF",X"FFFDFE",X"FFFEFD",X"FFFEFD",X"FFFDFF",X"FFFCFF",X"FFFBFF",X"FEFEFC",X"FFFFFD",X"FDFDFB",X"FFFFFD",X"FEFEFC",X"FDFDFD",X"FEFEFF",X"F4F2F5",X"3D342D",X"550700",X"B61E2B",X"C00B2C",X"C10E23",X"BF0E20",X"C00D2D",X"C21030",X"C31629",X"B01D25",X"8B0400",X"FFD9D8",X"FFFDFF",X"F5FFF7",X"F3FFFF",X"FBFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFCF9",X"FBFEED",X"CCE6CD",X"54953B",X"61B057",X"5CA44E",X"74AF5B",X"6DB053",X"67A753",X"6AA74A",X"66A344",X"68A152",X"76AB51",X"6A9345",X"CCE3C9",X"FBFFFA",X"FCFFF8",X"FEFFF4",X"FEFFF6",X"FEFFFA",X"FFFFFB",X"FFFFFA",X"FFFFF6",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FEFFFD",X"FDFFFC",X"FEFCFD",X"FFFCFF",X"FFFCFF",X"CBE1FF",X"0041A9",X"1673DD",X"0361D2",X"0772E4",X"0C79E0",X"0661D3",X"136CD2",X"0A6FE3",X"1B7DD6",X"0754B0",X"5D8DBE",X"F0FFFF",X"FBF4FF",X"FFFAFF",X"FBFFF3",X"FFFBFF",X"FFFAFF",X"FEF8FF",X"FEFCFF",X"FFFBF2",X"D1D076",X"D8D71A",X"DCCC1F",X"E0D40E",X"DBCD0C",X"E1D007",X"E4D100",X"E9D502",X"E6D30D",X"DFCF08",X"DFD400",X"E3DB1E",X"E3CF20",X"E7C853",X"9E855C",X"060000",X"0C0000",X"4D1106",X"67000B",X"AF040C",X"D60F14",X"ED040A",X"EF0007",X"DD081C",X"AA1229",X"4F0216",X"35212C",X"000A07",X"060002",X"110000",X"7B792C",X"B1B834",X"E6E241",X"DACE1A",X"D4CA06",X"DACB2A",X"969B47",X"000200",X"070016",X"00083F",X"1353AA",X"0C6ED3",X"0260C0",X"0B69CD",X"1C80EF",X"0052C6",X"1567D5",X"0858BB",X"3A5EB2",X"BCAAD2",X"BE9A8A",X"D87764",X"D86F52",X"D07A59",X"B08982",X"848BC1",X"335DC3",X"1264CA",X"057BC5",X"1067C4",X"226BC9",X"275FB2",X"29538D",X"26385E",X"241035",X"260024",X"5A0352",X"921C70",X"B11576",X"CF0E7B",X"C6016D",X"C10C6D",X"AF1064",X"9D1A5E",X"8D225A",X"4A1936",X"2D082A",X"070431",X"0C3875",X"165FAE",X"1A65C0",X"1865B5",X"1E6FB1",X"3669AB",X"14396D",X"0D1D37",X"150E16",X"34201F",X"635353",X"313237",X"0C1A25",X"0D2C2E",X"3A6367",X"317578",X"3EAFA9",X"019D88",X"00A286",X"01A283",X"12A185",X"0BB49D",X"19B59F",X"1F9D85",X"348370",X"012523",X"000B20",X"001647",X"225396",X"024097",X"B5DAFF"),
(X"FDFBFC",X"829593",X"0B7E61",X"26C4A3",X"00C29B",X"02C4A2",X"07BB9E",X"0ABD9F",X"00B79C",X"02D69B",X"32C2A9",X"357962",X"0F0004",X"19171A",X"B66B28",X"F48319",X"FF7000",X"FC7700",X"EE7800",X"FA8712",X"E57310",X"EA853D",X"D28B5F",X"502409",X"060000",X"000B0B",X"00211F",X"0E514A",X"136056",X"05564F",X"07585B",X"065863",X"096564",X"004F53",X"185D64",X"0B5558",X"005352",X"04605D",X"005655",X"126062",X"0B5554",X"144C4D",X"143033",X"11181E",X"00040A",X"000B09",X"001F14",X"006150",X"0FA0B3",X"23C5D4",X"1FDBE6",X"0BDAE2",X"00D4DF",X"04CFDE",X"10CEE4",X"14C9E4",X"00D7D9",X"05DCE1",X"00D4DF",X"00CDDC",X"00CCDC",X"06D5E5",X"05D7E6",X"07DBE7",X"02D7D1",X"03D3D3",X"06CFD6",X"10CAD7",X"1DC5D2",X"33C3CE",X"43BEC5",X"45B5B7",X"487570",X"001310",X"000100",X"110907",X"030000",X"000800",X"284D21",X"609358",X"79A165",X"8DB775",X"77AA5F",X"7EBB6B",X"6FB05E",X"7BB666",X"82B163",X"93B568",X"7BA86F",X"1A2014",X"060010",X"7F1150",X"DF177A",X"E01080",X"B70166",X"E076B8",X"FFE7F6",X"FFFCFF",X"F9FFFF",X"FFFEFF",X"FFF9FB",X"FEFFFF",X"FCFEFD",X"FFFDFF",X"FFF9FF",X"E5F0EC",X"498271",X"006F53",X"1EBEA2",X"0BCCAD",X"00AE96",X"0FB59F",X"0FD0B1",X"03B49A",X"07B59A",X"16AE97",X"3FC8AE",X"D5F7F8",X"FEF9FF",X"F9FFFD",X"FFFAFF",X"FFFCFF",X"FFFDFE",X"FFFEFD",X"FFFEFD",X"FFFDFF",X"FFFCFF",X"FFFBFF",X"FEFEFC",X"FFFFFD",X"FDFDFB",X"FFFFFD",X"FEFEFC",X"FDFDFD",X"FEFEFF",X"F4F2F5",X"3C332C",X"530500",X"B41C29",X"BD0829",X"BD0A1F",X"BB0A1C",X"BE0B2B",X"BF0D2D",X"BD1023",X"AE1B23",X"8B0400",X"FED8D7",X"FFFDFF",X"F6FFF8",X"F4FFFF",X"FBFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FCFBFF",X"FDF9F6",X"FFFFF1",X"CDE7CE",X"55963C",X"61B057",X"5DA54F",X"68A34F",X"70B356",X"6CAC58",X"7EBB5E",X"5F9C3D",X"629B4C",X"73A84E",X"719A4C",X"C9E0C6",X"FBFFFA",X"FCFFF8",X"FEFFF4",X"FEFFF6",X"FEFFFA",X"FFFFFB",X"FFFFFA",X"FFFFF6",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FEFFFD",X"FDFFFC",X"FEFCFD",X"FFFCFF",X"FFFCFF",X"BCD2FF",X"084BB3",X"1774DE",X"0664D5",X"0974E6",X"0F7CE3",X"0D68DA",X"116AD0",X"0368DC",X"0668C1",X"0C59B5",X"6A9ACB",X"EBFCFF",X"FFFBFF",X"F8F3F9",X"FBFFF3",X"FDF8FF",X"FFFAFF",X"FFFAFF",X"FFFEFF",X"FFFFF6",X"DEDD83",X"D6D518",X"DACA1D",X"D8CC06",X"E6D817",X"E4D30A",X"DAC700",X"E7D300",X"DDCA04",X"E6D60F",X"DCD100",X"E4DC1F",X"EBD728",X"A98A15",X"170000",X"272016",X"120500",X"5F2318",X"96273A",X"C41921",X"CE070C",X"ED040A",X"E80000",X"D20011",X"B11930",X"520519",X"2D1924",X"172724",X"060002",X"867563",X"DAD88B",X"DAE15D",X"C9C524",X"D4C814",X"E1D713",X"D9CA29",X"2A2F00",X"000200",X"241733",X"2E376E",X"2969C0",X"1C7EE3",X"005ABA",X"0664C8",X"005ECD",X"136CE0",X"1264D2",X"0050B3",X"1F4397",X"6B5981",X"A88474",X"D97865",X"DF7659",X"DE8867",X"966F68",X"282F65",X"4B75DB",X"0F61C7",X"1288D2",X"1970CD",X"2871CF",X"043C8F",X"001953",X"001238",X"3A264B",X"4E114C",X"7B2473",X"911B6F",X"B01475",X"D00F7C",X"C6016D",X"B80364",X"AC0D61",X"8B084C",X"60002D",X"1F000B",X"160013",X"2A2754",X"36629F",X"2770BF",X"115CB7",X"1D6ABA",X"1364A6",X"093C7E",X"000A3E",X"00051F",X"0B040C",X"685453",X"7A6A6A",X"65666B",X"1E2C37",X"001F21",X"00171B",X"002528",X"14857F",X"19B5A0",X"03B094",X"0DAE8F",X"0D9C80",X"009C85",X"0EAA94",X"18967E",X"004532",X"052927",X"001227",X"1D3D6E",X"4273B6",X"08469D",X"BBE0FF"),
(X"FFFFFF",X"998D91",X"095842",X"34C4A3",X"00C39A",X"00C2A1",X"06C1A2",X"0DC2A1",X"09BFA9",X"1AC6AE",X"31C8A7",X"355A52",X"0B010A",X"592B11",X"E67E25",X"FF7C0F",X"F98000",X"FF8009",X"F86A00",X"FF7209",X"FF8317",X"F37F10",X"F5861D",X"E0740F",X"6F2700",X"240000",X"160F09",X"011A21",X"1F4B54",X"205D60",X"07524E",X"045954",X"036163",X"00585D",X"086167",X"065D64",X"005359",X"0D5E61",X"116361",X"045650",X"155756",X"084C4D",X"195C62",X"205B63",X"00242D",X"00111B",X"00090D",X"000104",X"010012",X"334F5B",X"50979B",X"4EC2C1",X"33CCC9",X"16C9C6",X"0AD2CF",X"00D2CE",X"13D5DE",X"0CD7DD",X"01D6DA",X"00D1D4",X"05D6DA",X"08D3D7",X"08D2D2",X"09D1CE",X"07D9EA",X"01D7E2",X"01DCE0",X"03E2E1",X"01D8DA",X"03CFDA",X"0DCBE3",X"15C9EA",X"29CFE5",X"0FA3AF",X"1E9494",X"045B53",X"00120B",X"000E0C",X"000105",X"060004",X"394231",X"6B8265",X"83AA7B",X"8FBA82",X"8AB276",X"83AD6B",X"7FB569",X"6FB55F",X"75A969",X"28291B",X"08000D",X"622044",X"AF1A5A",X"E5247F",X"CF066E",X"DF4198",X"FFDAED",X"FFFAFF",X"FAFFFF",X"FFFFFF",X"FFFAFC",X"FCFEFD",X"FAFEFD",X"FFFEFF",X"EBFFFF",X"FFFCFF",X"888D87",X"000104",X"4EAB99",X"4CAEA1",X"15AC89",X"2BBC93",X"15B496",X"17C7A3",X"00C196",X"12B795",X"00B98A",X"B8F4E8",X"FBFFFE",X"F8FAF5",X"FCFDFF",X"FDFEFF",X"FDFEFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FEFEFC",X"FFFFFD",X"FDFDFB",X"FFFFFF",X"FEFEFE",X"FDFDFD",X"FEFEFE",X"F3F3F3",X"30393E",X"530505",X"C11432",X"D00037",X"CB0030",X"C80128",X"CE012A",X"D40320",X"E2002D",X"D20B32",X"AB0012",X"FFD2E9",X"FEFBFF",X"FBFFFE",X"F6FFFF",X"FEFFF9",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFCFF",X"FFF9F9",X"FEFFF1",X"C7DEC4",X"5F953D",X"6BAF58",X"65A952",X"609E49",X"6BA05A",X"71A368",X"72A362",X"72A361",X"7BAA74",X"79A276",X"75936D",X"CBDFC4",X"FFFCFF",X"FFFDFF",X"FFFEFF",X"FFFDFF",X"FFFCFF",X"FFFBFF",X"FFFCFF",X"FFFDFF",X"FCFFFB",X"FCFFFB",X"FCFFFB",X"FCFFFB",X"FDFFFC",X"FEFCFD",X"FFFCFF",X"FFFCFF",X"C0D4F7",X"0A4CC6",X"1270E4",X"1266E2",X"0F70E5",X"006DCC",X"0362D8",X"0E6EC2",X"185DA8",X"3A74B3",X"24478B",X"7488A1",X"E9F3EB",X"F8F7FD",X"FFFEFF",X"FCFBF9",X"FFFAFE",X"FFFFEE",X"FFFCFF",X"FDFCFF",X"FFFFF3",X"E9E987",X"D0D300",X"D8C90A",X"D8CF06",X"E8DC14",X"D1C300",X"E5D50C",X"DAD100",X"E2DF00",X"D4D110",X"D9D33D",X"CCCC54",X"8A8F4C",X"000700",X"0F161E",X"0C0009",X"4C0515",X"B40E24",X"F9061C",X"D90106",X"D6050A",X"D50000",X"EF0609",X"EA0406",X"D7050E",X"A10D1D",X"46000C",X"171103",X"0A000B",X"767062",X"CDD069",X"C1C816",X"D5D10E",X"DFC607",X"EEC400",X"D4C029",X"716501",X"0A0200",X"271F2C",X"2A3867",X"2358A6",X"1265CD",X"0261D5",X"0F6BD0",X"086ACF",X"1067D1",X"0D63D2",X"1071E2",X"166ADE",X"0A49B2",X"004092",X"325CB2",X"3B6AB0",X"2662AA",X"0051AD",X"035EC7",X"166ED0",X"276FC3",X"2967B2",X"215168",X"1C2C4E",X"26103E",X"27002A",X"500038",X"8E0058",X"BC0B73",X"C20772",X"C9006B",X"DC0676",X"C40063",X"B01769",X"9D2F6C",X"6C2148",X"1F0010",X"1B2622",X"083329",X"0F181F",X"121734",X"285B92",X"1263B2",X"296BBF",X"214A82",X"072740",X"080812",X"0C0807",X"2B1D10",X"866A54",X"997255",X"986F51",X"99775B",X"856A4D",X"190000",X"0A0000",X"1C2124",X"142C30",X"386369",X"3A8483",X"2B998E",X"1EA692",X"2CADA8",X"3D988F",X"16453F",X"051B29",X"152F60",X"003080",X"0757B6",X"0C6ED1",X"0035A7",X"B5D3FF"),
(X"FEFEFE",X"978B8F",X"003D27",X"2EBE9D",X"00BD94",X"00BE9D",X"05C0A1",X"07BC9B",X"06BCA6",X"16C2AA",X"1CB392",X"00231B",X"060005",X"73452B",X"F48C33",X"F67205",X"FB8200",X"FF7A03",X"FF8012",X"FC6D04",X"FC790D",X"ED790A",X"E3740B",X"FE922D",X"BF7747",X"3A0D00",X"0C0500",X"00141B",X"00151E",X"155255",X"0B5652",X"156A65",X"005D5F",X"005C61",X"005359",X"085F66",X"0B5E64",X"0B5C5F",X"166866",X"00524C",X"034544",X"105455",X"0E5157",X"09444C",X"27525B",X"1C343E",X"071216",X"050A0D",X"020113",X"000713",X"00171B",X"006665",X"1EB7B4",X"27DAD7",X"1BE3E0",X"03D8D4",X"0BCDD6",X"05D0D6",X"04D9DD",X"01D8DB",X"08D9DD",X"00CBCF",X"06D0D0",X"12DAD7",X"02D4E5",X"00D0DB",X"00D5D9",X"00DFDE",X"03DADC",X"06D2DD",X"0ECCE4",X"16CAEB",X"1CC2D8",X"31C5D1",X"4EC4C4",X"449B93",X"2D665F",X"2C4947",X"04090D",X"080006",X"000500",X"000A00",X"163D0E",X"406B33",X"6F975B",X"7FA967",X"7FB569",X"87CD77",X"84B878",X"2B2C1E",X"06000B",X"310013",X"950040",X"CF0E69",X"DA1179",X"AE1067",X"F5CEE1",X"FFF7FF",X"F8FEFE",X"FFFFFF",X"FFFCFE",X"FEFFFF",X"FAFEFD",X"FEFCFD",X"EEFFFF",X"FFFCFF",X"7D827C",X"000306",X"005B49",X"2E9083",X"10A784",X"25B68D",X"24C3A5",X"1ACAA6",X"00BA8F",X"23C8A6",X"02BC8D",X"A7E3D7",X"FBFFFE",X"FEFFFB",X"FCFDFF",X"FDFEFF",X"FDFEFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FEFEFC",X"FFFFFD",X"FDFDFB",X"FFFFFF",X"FEFEFE",X"FDFDFD",X"FEFEFE",X"F3F3F3",X"30393E",X"530505",X"C11432",X"CF0036",X"CB0030",X"C70027",X"CC0028",X"D1001D",X"E0002B",X"D30C33",X"AD0014",X"FFD1E8",X"FCF9FF",X"FBFFFE",X"F7FFFF",X"FEFFF9",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FBF5FF",X"FFF9F9",X"FEFFF1",X"CBE2C8",X"669C44",X"6DB15A",X"6DB15A",X"77B560",X"72A761",X"79AB70",X"72A362",X"6B9C5A",X"54834D",X"3B6438",X"001300",X"ABBFA4",X"FFFCFF",X"FFFDFF",X"FFFEFF",X"FFFDFF",X"FFFCFF",X"FFFBFF",X"FFFCFF",X"FFFDFF",X"FCFFFB",X"FCFFFB",X"FCFFFB",X"FCFFFB",X"FDFFFC",X"FEFCFD",X"FFFCFF",X"FFFCFF",X"CDE1FF",X"0F51CB",X"1573E7",X"1064E0",X"0B6CE1",X"006BCA",X"0D6CE2",X"1272C6",X"2166B1",X"1E5897",X"000347",X"354962",X"E4EEE6",X"FFFEFF",X"FBF9FA",X"FEFDFB",X"FFFDFF",X"FFFFEF",X"FDFAFF",X"FBFAFF",X"FFFDF1",X"F2F290",X"CED100",X"E1D213",X"D6CD04",X"D5C901",X"E0D20D",X"E7D70E",X"DDD400",X"D5D200",X"D7D413",X"E3DD47",X"85850D",X"070C00",X"192112",X"10171F",X"1E111B",X"641D2D",X"BA142A",X"EF0012",X"D80005",X"D10005",X"DC0107",X"E90003",X"E30000",X"DD0B14",X"AE1A2A",X"621A28",X"120C00",X"261C27",X"080200",X"4E5100",X"C7CE1C",X"E3DF1C",X"D4BB00",X"EEC400",X"DDC932",X"D2C662",X"3C3410",X"040009",X"000231",X"0E4391",X"1467CF",X"0463D7",X"0561C6",X"1072D7",X"0158C2",X"0C62D1",X"0465D6",X"0559CD",X"2160C9",X"1E66B8",X"204AA0",X"16458B",X"2561A9",X"1667C3",X"0F6AD3",X"146CCE",X"2169BD",X"013F8A",X"00162D",X"000123",X"2E1846",X"59245C",X"83236B",X"A1106B",X"C7167E",X"C20772",X"CF0571",X"CC0066",X"D30A72",X"AA1163",X"841653",X"3F001B",X"1A000B",X"1A2521",X"164137",X"141D24",X"00001B",X"002A61",X"0F60AF",X"1254A8",X"00225A",X"000922",X"000009",X"676362",X"8D7F72",X"A0846E",X"9F785B",X"AB8264",X"A58367",X"816649",X"7D6062",X"6D5F5F",X"23282B",X"152D31",X"000C12",X"004544",X"00695E",X"08907C",X"33B4AF",X"2C877E",X"001610",X"0F2533",X"051F50",X"2C61B1",X"1363C2",X"1072D5",X"053AAC",X"BBD9FF"),
(X"FAFFFE",X"9F8A8F",X"00331B",X"2BBB97",X"00BB94",X"04BFA2",X"0CC7AA",X"00BE99",X"03B39F",X"34B8AB",X"18765E",X"0C000B",X"0C0100",X"BC641A",X"F8841D",X"FF790F",X"FC7C11",X"F47B0A",X"FD860E",X"F77A00",X"FF7300",X"FF7200",X"FF7C09",X"F67C0D",X"F88417",X"C76615",X"561200",X"220000",X"1F0700",X"050300",X"20382A",X"194538",X"196460",X"055C56",X"005652",X"005D5D",X"0B5C60",X"095356",X"095553",X"0E605A",X"135F55",X"06534D",X"0A5457",X"10545F",X"1B5666",X"0D4755",X"0C4B52",X"064A4D",X"002A17",X"002A1C",X"00130C",X"00070A",X"011A21",X"1B4E51",X"409B96",X"52CCBF",X"3ECED9",X"2FD2DB",X"1FD8DD",X"0CD3DA",X"0FDAE1",X"06CFD9",X"05CED8",X"01CDD4",X"0DE1E4",X"09D8E0",X"09D2E2",X"0ED1E7",X"0CCFE5",X"0BD0E3",X"0BD5E3",X"06D5DD",X"0DD7EB",X"06D1DF",X"04D3D9",X"07D4D7",X"0FD1D0",X"1AC5BF",X"008A7E",X"005243",X"000F10",X"000C0C",X"000200",X"010100",X"000600",X"384B37",X"50684E",X"6C8366",X"7F9580",X"38302E",X"000600",X"0C1500",X"380E0F",X"86264C",X"CB2571",X"D2005B",X"F6C6DC",X"FFF8FF",X"F8FCFD",X"FDFDFD",X"FFFDFF",X"FEFFFF",X"FBFFFF",X"FBFDFC",X"FBF9FF",X"FCFCF2",X"B2BC9A",X"1A0600",X"220C00",X"010000",X"16221E",X"18362C",X"5A7481",X"498689",X"3EA39D",X"459F9D",X"259A8A",X"B1DADE",X"FBFFFF",X"FAF7FF",X"F7FFFD",X"FAFFFE",X"FAFFFF",X"FBFFFF",X"FBFFFF",X"FBFFFF",X"FBFFFF",X"FBFFFD",X"FFFDFE",X"FFFEFF",X"FEFCFF",X"FFFEFF",X"FFFDFF",X"FDFDFD",X"FEFEFE",X"F3F3F3",X"373334",X"510200",X"B9152D",X"C50030",X"C50328",X"C4011F",X"CA001F",X"CD0016",X"C60611",X"BF161B",X"A50000",X"FFD5D6",X"FBFAFF",X"FFFCF9",X"FFFEFF",X"FFFAFD",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFDFF",X"FFFEFF",X"FBFEF5",X"D1DAD5",X"7E925F",X"859D7B",X"6C896D",X"6E8C74",X"76796E",X"53544F",X"353537",X"3A3F3B",X"000107",X"07052A",X"080021",X"CAC0BF",X"F8FFFF",X"F9FFFD",X"F9FFFB",X"F9FFFD",X"F9FFFF",X"F9FFFF",X"F9FFFF",X"F9FFFB",X"FEFFFB",X"FEFFFD",X"FFFFFD",X"FFFFFF",X"FFFDFE",X"FEFCFD",X"FEFEFE",X"FFFFFF",X"C6E1F4",X"075AC4",X"0B7BEB",X"0164C9",X"0A6CC7",X"1B74C8",X"2E65CA",X"1D458D",X"0B2639",X"00040D",X"261C1A",X"080300",X"CBCEB3",X"F6FAFF",X"F8F8FF",X"FFF8FF",X"FFFCFF",X"FEFEF2",X"FBF6FF",X"FDFCFF",X"FFFFF3",X"F9F4B2",X"D5D213",X"E9DE0A",X"E4CB00",X"E8CF01",X"E3CB07",X"D2BC07",X"DFCF24",X"EBE249",X"CEC75C",X"6B6124",X"000100",X"002319",X"004D41",X"0A4847",X"1B1716",X"5D0803",X"D2222D",X"EB001B",X"D30207",X"D40C0F",X"DB080E",X"DB0409",X"D70707",X"DB080F",X"CB111C",X"931719",X"483141",X"0A1B13",X"031F13",X"030000",X"9B8755",X"E9E462",X"CCD01B",X"D9D619",X"DBCD00",X"F8D814",X"C9AB29",X"0B0500",X"000301",X"0F1A30",X"2C4C87",X"2064C5",X"0D5DCC",X"0A67C6",X"1069CF",X"0C69E2",X"0A6FE3",X"0D63CA",X"1762C8",X"0264CF",X"1C67CD",X"0C5FBB",X"246AC0",X"3E6CBA",X"3C5D92",X"36516E",X"1A163B",X"1F0034",X"2F001F",X"6E0442",X"960955",X"BC1B78",X"CA1282",X"DA0A82",X"C80066",X"C80C63",X"C00F60",X"B01E65",X"87295D",X"3B0D2A",X"070005",X"061A11",X"073F22",X"0E6135",X"335F3B",X"114D34",X"001419",X"000A2D",X"26254F",X"09122F",X"000213",X"2F1B27",X"8B7665",X"8F7D69",X"8E7E67",X"8F7A5F",X"8F7051",X"A57F58",X"AA8153",X"8B632F",X"977665",X"AC8F7F",X"826B5B",X"130500",X"0A0600",X"000100",X"010C10",X"24353C",X"3A565A",X"081319",X"060C1C",X"00173F",X"1C5CA3",X"136AC9",X"1867D0",X"2C69D4",X"0342A1",X"BCDDFF"),
(X"FBFFFF",X"A18C91",X"003D25",X"2CBC98",X"01C19A",X"0CC7AA",X"14CFB2",X"03C39E",X"10C0AC",X"2AAEA1",X"004C34",X"0B000A",X"382D17",X"DC843A",X"EF7B14",X"FF780E",X"FC7C11",X"F77E0D",X"F37C04",X"FB7E00",X"FF7F03",X"FF7200",X"FA7401",X"F97F10",X"F17D10",X"E38231",X"CF8B5C",X"835641",X"180000",X"030100",X"000900",X"002B1E",X"0D5854",X"156C66",X"046460",X"026060",X"0A5B5F",X"065053",X"0E5A58",X"0A5C56",X"065248",X"08554F",X"054F52",X"125661",X"0E4959",X"134D5B",X"16555C",X"165A5D",X"235C49",X"0E3E30",X"02231C",X"011619",X"000C13",X"000F12",X"00322D",X"006B5E",X"1FAFBA",X"26C9D2",X"20D9DE",X"0CD3DA",X"09D4DB",X"0CD5DF",X"0ED7E1",X"08D4DB",X"00CED1",X"00CFD7",X"09D2E2",X"11D4EA",X"0FD2E8",X"10D5E8",X"0DD7E5",X"05D4DC",X"12DCF0",X"07D2E0",X"01D0D6",X"0BD8DB",X"11D3D2",X"1EC9C3",X"3CCABE",X"44BDAE",X"4E8081",X"2A4848",X"000501",X"060600",X"000500",X"000800",X"000C00",X"000B00",X"162C17",X"19110F",X"000E03",X"000800",X"1E0000",X"500016",X"CB2571",X"CB0054",X"F5C5DB",X"FFF9FF",X"F8FCFD",X"FBFBFB",X"FFFBFD",X"FDFFFE",X"FBFFFF",X"FCFEFD",X"FCFAFF",X"FFFFF6",X"BFC9A7",X"57432A",X"160000",X"1C1B16",X"000602",X"001309",X"000613",X"001316",X"00544E",X"1C7674",X"087D6D",X"AFD8DC",X"F6FAFF",X"FFFDFF",X"F7FFFD",X"FAFFFE",X"FAFFFF",X"FBFFFF",X"FBFFFF",X"FBFFFF",X"FBFFFF",X"FBFFFD",X"FFFDFE",X"FFFEFF",X"FEFCFF",X"FFFEFF",X"FFFDFF",X"FDFDFD",X"FEFEFE",X"F3F3F3",X"3A3637",X"540500",X"BB172F",X"C70132",X"C8062B",X"C80523",X"CE0223",X"D1031A",X"CC0C17",X"C1181D",X"A60000",X"FFD7D8",X"FDFCFF",X"FFFCF9",X"FFFEFF",X"FFFAFD",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFAFF",X"FCFAFB",X"FAFDF4",X"D9E2DD",X"5F7340",X"4B6341",X"09260A",X"000F00",X"080B00",X"000100",X"020204",X"000200",X"000309",X"232146",X"03001C",X"C8BEBD",X"F8FFFF",X"F9FFFD",X"F9FFFB",X"F9FFFD",X"F9FFFF",X"F9FFFF",X"F9FFFF",X"F9FFFB",X"FEFFFB",X"FEFFFD",X"FFFFFD",X"FFFFFF",X"FFFDFE",X"FEFCFD",X"FEFEFE",X"FFFFFF",X"CAE5F8",X"1669D3",X"0474E4",X"0C6FD4",X"0F71CC",X"0E67BB",X"063DA2",X"000E56",X"00182B",X"00020B",X"080000",X"423D15",X"D4D7BC",X"F8FCFF",X"FEFEFF",X"FDF1FF",X"FFFBFF",X"FDFDF1",X"FDF8FF",X"FFFEFF",X"FFFFF4",X"FBF6B4",X"D7D415",X"E1D602",X"E7CE00",X"F2D90B",X"E0C804",X"F0DA25",X"E2D227",X"C4BB22",X"898217",X"0E0400",X"010504",X"4E8379",X"459D91",X"2F6D6C",X"080403",X"550000",X"BE0E19",X"EC001C",X"CF0003",X"DC1417",X"D40107",X"DF080D",X"E41414",X"D6030A",X"CD131E",X"8B0F11",X"2B1424",X"33443C",X"122E22",X"15120B",X"140000",X"868100",X"E6EA35",X"D1CE11",X"DED000",X"DABA00",X"F9DB59",X"958F5B",X"000200",X"172238",X"001954",X"1B5FC0",X"0F5FCE",X"0663C2",X"116AD0",X"0055CE",X"0469DD",X"0B61C8",X"206BD1",X"0769D4",X"0F5AC0",X"1B6ECA",X"1D63B9",X"1D4B99",X"08295E",X"000522",X"09052A",X"300145",X"641E54",X"922866",X"A51864",X"B41370",X"C00878",X"D10179",X"CE006C",X"CA0E65",X"C11061",X"A31158",X"610337",X"1E000D",X"10040E",X"2D4138",X"225A3D",X"2B7E52",X"2A5632",X"27634A",X"033439",X"021033",X"000026",X"000623",X"16192A",X"533F4B",X"988372",X"73614D",X"6A5A43",X"897459",X"6D4E2F",X"9B754E",X"976E40",X"A37B47",X"927160",X"775A4A",X"9C8575",X"6F6154",X"363229",X"2D3130",X"000307",X"00050C",X"00080C",X"00080E",X"010717",X"1D3961",X"2B6BB2",X"1B72D1",X"1362CB",X"2562CD",X"0241A0",X"BBDCFF"),
(X"F6FFFD",X"9B888A",X"004B2E",X"25BC93",X"04BE99",X"10BCA6",X"0FC7AB",X"00C39B",X"24C7B2",X"11946C",X"0D0B0E",X"0A0002",X"885424",X"E69520",X"FC7701",X"F27207",X"F78501",X"F58205",X"FE8711",X"FC800E",X"F57301",X"FF790A",X"FB7409",X"FE7610",X"FF7F02",X"F97C06",X"F28619",X"E98925",X"C26B1B",X"763300",X"310900",X"0D000B",X"201F1D",X"304341",X"225350",X"165E5D",X"095D5F",X"035D5E",X"086665",X"005654",X"00525B",X"086366",X"005D57",X"025F54",X"01584F",X"0A5F58",X"095E5B",X"005556",X"08555F",X"125F67",X"1B6067",X"083A41",X"052029",X"0C1620",X"00030C",X"000309",X"000A0A",X"234A47",X"448F8B",X"4CBABB",X"3FC9CC",X"2CCFD6",X"14CFD4",X"07D4D7",X"0FD3E3",X"0BD1DE",X"09D3DD",X"06D7DB",X"02D6D7",X"01D9D8",X"02DAD9",X"00D6D5",X"00CFD1",X"06DADB",X"02D4D5",X"06D5DB",X"07D5E3",X"06CFE3",X"0DCDE4",X"0EC8DD",X"1DD2E7",X"1AC7D5",X"19B2B8",X"108992",X"004858",X"000E23",X"00091E",X"000C1C",X"000716",X"0A0A12",X"030700",X"483912",X"2D1800",X"000100",X"5E3148",X"8D0E3B",X"EEBAD1",X"FFF8FF",X"F8FCFD",X"FBFBFB",X"FFFCFD",X"FCFEFD",X"FBFFFF",X"FAFEFD",X"F9F9FF",X"FFFAEC",X"DEEAA8",X"CB975D",X"1A0600",X"081700",X"14070E",X"3B1934",X"4E0E28",X"2C0011",X"18000B",X"1B000C",X"190010",X"98788D",X"FFF4FE",X"FFF9FC",X"FFFCF9",X"FFFCFC",X"FFFCFF",X"FFFCFF",X"FFFCFF",X"FFFDFF",X"FFFEFB",X"FFFFFA",X"FFFDFF",X"FFFEFF",X"FEFCFF",X"FFFEFF",X"FFFDFF",X"FDFDFD",X"FEFEFE",X"F3F3F1",X"39363F",X"470A09",X"A02132",X"A71031",X"AC1325",X"B21123",X"B80E32",X"B80F36",X"BA132F",X"B21A2F",X"9D0009",X"FFDBDD",X"FBFFFF",X"FFFFF7",X"F5FFFF",X"FDFFFA",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFF9FC",X"FEFEFE",X"F8FEFE",X"C2C7DA",X"020901",X"00081D",X"000127",X"000332",X"000D3F",X"00275D",X"003476",X"003975",X"0F4E91",X"184EBB",X"0B3CA5",X"A4DAFE",X"FFFAFF",X"FFFDFF",X"FFFDFD",X"FFFDFD",X"FFFDFF",X"FFFDFF",X"FFFDFF",X"FFFEFD",X"FFFEFF",X"FFFDFF",X"FFFDFF",X"FFFCFF",X"FFFCFF",X"FDFDFD",X"FBFFFA",X"FBFFFA",X"EEFBF4",X"548ED7",X"1854B4",X"3D5A92",X"334865",X"1C2E42",X"0A0F12",X"040300",X"040900",X"4E3F00",X"BDA123",X"D3C530",X"ECF19F",X"F8FFF6",X"F4F8E9",X"FFF7FA",X"FDFFFA",X"FFFFEC",X"FFFCFF",X"FDFCF8",X"FFFEFB",X"FFF0E3",X"E1D44A",X"D8C705",X"E4DB1E",X"DDD326",X"E5DB46",X"CBC555",X"747239",X"000100",X"00030B",X"000F07",X"004428",X"29B38F",X"36CEA5",X"08704F",X"000800",X"531113",X"A6120E",X"E41706",X"E8090C",X"D8000C",X"ED001A",X"E3000B",X"E4030B",X"EA0710",X"CF0417",X"9C1420",X"160B13",X"21635F",X"2D9E82",X"003B1A",X"000E09",X"080206",X"988F54",X"E7D648",X"D0C921",X"E6DD28",X"C4BE10",X"D3D351",X"736F30",X"040000",X"1A213B",X"173058",X"335AB7",X"106DCD",X"005AC6",X"0957C6",X"176AD0",X"0059B9",X"0C5CBB",X"1862BB",X"2360A3",X"375B97",X"232E5C",X"01001B",X"1E001A",X"520030",X"6F003D",X"A1156C",X"BF1487",X"C50073",X"D80072",X"CF006D",X"D50D7A",X"C50670",X"C2237F",X"961E66",X"6C1F3F",X"2C000D",X"361424",X"12060A",X"2D493A",X"0F5934",X"116D3A",X"075A26",X"0D7236",X"116A32",X"104821",X"010E07",X"292033",X"281D2E",X"281D1B",X"0F0000",X"1C0000",X"160000",X"100000",X"0B0000",X"0C0000",X"261815",X"342B22",X"847E72",X"8D715B",X"947259",X"8B6349",X"A88066",X"89674E",X"947B67",X"504031",X"0A0000",X"0B0000",X"25241F",X"0B191C",X"16263D",X"1C2F5A",X"345491",X"3369B1",X"226CB7",X"064894",X"C2E4FF"),
(X"F8FFFF",X"9B888A",X"08583B",X"28BF96",X"07C19C",X"0DB9A3",X"0BC3A7",X"00C49C",X"25C8B3",X"04875F",X"030104",X"0A0002",X"9D6939",X"EE9D28",X"FF850F",X"FF8116",X"FA8804",X"FF9114",X"F27B05",X"FD810F",X"FF800E",X"F97304",X"F36C01",X"FF7A14",X"FE7400",X"FE810B",X"F28619",X"E3831F",X"E99242",X"D79460",X"593127",X"0D000B",X"0F0E0C",X"000604",X"0F403D",X"0F5756",X"065A5C",X"0B6566",X"005453",X"005D5B",X"085F68",X"005659",X"005C56",X"036055",X"045B52",X"00544D",X"116663",X"01595A",X"0F5C66",X"004C54",X"13585F",X"23555C",X"314C55",X"2A343E",X"050E17",X"061319",X"000C0C",X"000C09",X"001814",X"005253",X"079194",X"1FC2C9",X"17D2D7",X"13E0E3",X"14D8E8",X"07CDDA",X"00C9D3",X"00D1D5",X"02D6D7",X"04DCDB",X"05DDDC",X"01D9D8",X"05DCDE",X"02D6D7",X"00D1D2",X"0CDBE1",X"03D1DF",X"05CEE2",X"0BCBE2",X"14CEE3",X"14C9DE",X"16C3D1",X"30C9CF",X"4EC7D0",X"4A9DAD",X"52899E",X"3C6277",X"395D6D",X"233D4C",X"010109",X"050900",X"AE9F78",X"A99477",X"050600",X"33061D",X"730021",X"E1ADC4",X"FFF5FF",X"F8FCFD",X"FDFDFD",X"FFFEFF",X"FCFEFD",X"FBFFFF",X"F9FDFC",X"FBFBFF",X"FFFAEC",X"F2FEBC",X"EDB97F",X"A5915C",X"000B00",X"0C0006",X"4F2D48",X"874761",X"57263C",X"3C162F",X"390E2A",X"321029",X"321227",X"F6E5EF",X"FFFAFD",X"FFFCF9",X"FFFCFC",X"FFFCFF",X"FFFCFF",X"FFFCFF",X"FFFDFF",X"FFFEFB",X"FFFFFA",X"FFFDFF",X"FFFEFF",X"FEFCFF",X"FFFEFF",X"FFFDFF",X"FDFDFD",X"FEFEFE",X"F3F3F1",X"333039",X"400302",X"98192A",X"9E0728",X"A40B1D",X"AC0B1D",X"B2082C",X"B30A31",X"B10A26",X"A81025",X"960002",X"FCD8DA",X"FBFFFF",X"FFFFF7",X"F6FFFF",X"FEFFFB",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFCFF",X"FCFCFC",X"FBFFFF",X"CBD0E3",X"000300",X"1B2338",X"293B61",X"34507F",X"265B8D",X"295E94",X"2C61A3",X"2F6AA6",X"3473B6",X"2D63D0",X"194AB3",X"9FD5F9",X"FFFAFF",X"FFFDFF",X"FFFDFD",X"FFFDFD",X"FFFDFF",X"FFFDFF",X"FFFDFF",X"FFFEFD",X"FFFEFF",X"FFFDFF",X"FFFDFF",X"FFFCFF",X"FFFCFF",X"FDFDFD",X"FBFFFA",X"FBFFFA",X"F5FFFB",X"75AFF8",X"003696",X"112E66",X"000B28",X"000317",X"000205",X"1E1D01",X"888D4D",X"D2C368",X"FBDF61",X"D4C631",X"DDE290",X"F6FFF4",X"FEFFF3",X"FFF6F9",X"FBFDF8",X"FFFFEC",X"FFFCFF",X"FBFAF6",X"FFFEFB",X"FFFAED",X"F1E45A",X"DBCA08",X"E0D71A",X"E0D629",X"C5BB26",X"686200",X"0D0B00",X"0C0E09",X"1A272F",X"5D746C",X"4EB296",X"2AB490",X"24BC93",X"40A887",X"001308",X"400000",X"A6120E",X"DB0E00",X"E10205",X"D8000C",X"EC0019",X"F2031A",X"EA0911",X"E10007",X"D3081B",X"910915",X"0C0109",X"0D4F4B",X"59CAAE",X"3D8766",X"000702",X"050003",X"0E0500",X"BDAC1E",X"E6DF37",X"D8CF1A",X"DDD729",X"D1D14F",X"938F50",X"060100",X"080F29",X"00153D",X"052C89",X"1B78D8",X"0B71DD",X"1C6AD9",X"1265CB",X"1C79D9",X"1767C6",X"347ED7",X"205DA0",X"000440",X"000634",X"090223",X"340F30",X"772555",X"A0276E",X"AC2077",X"B60B7E",X"CC057A",X"D4006E",X"CD006B",X"D60E7B",X"C70872",X"A80965",X"700040",X"3A000D",X"370018",X"310F1F",X"100408",X"254132",X"226C47",X"076330",X"136632",X"006529",X"1A733B",X"1C542D",X"0E1B14",X"170E21",X"120718",X"261B19",X"3C2A16",X"512A23",X"3B1C17",X"503B36",X"342522",X"0D0000",X"0C0000",X"070000",X"060000",X"4B2F19",X"704E35",X"8C644A",X"997157",X"B49279",X"846B57",X"8A7A6B",X"6F6259",X"584A41",X"010000",X"000407",X"000219",X"000934",X"12326F",X"00337B",X"09539E",X"00327E",X"B4D6F9"),
(X"FFFAFF",X"839B9B",X"00785C",X"30C9AD",X"10B799",X"09BC9C",X"0AC9AA",X"16C6B1",X"4AAC9D",X"194949",X"030002",X"523525",X"C2956C",X"CB8758",X"D17F59",X"D18063",X"C77952",X"C68754",X"D8924D",X"EF8A38",X"F48029",X"EB7921",X"EA7410",X"FC7A02",X"F86D06",X"FC7A0A",X"F88005",X"EE7B00",X"FB830B",X"F97F1C",X"E07726",X"7A2800",X"190000",X"150000",X"140502",X"0F1316",X"223E41",X"2E6260",X"145F5A",X"00534E",X"04554F",X"085A58",X"035256",X"0F5D5F",X"095354",X"0C5B58",X"0D6362",X"005E5E",X"125659",X"125B62",X"03525F",X"0A606F",X"035968",X"13666E",X"095555",X"054E47",X"002C2B",X"002629",X"001219",X"00030A",X"000205",X"0D201E",X"335E57",X"4D8A83",X"4FBECF",X"4ECAD6",X"34C3CB",X"22C7CB",X"14CDD0",X"06D0D4",X"08D9E0",X"00D4DE",X"00D3D5",X"08DCDF",X"06D6DA",X"03CED2",X"0CD7DB",X"03D1D1",X"05D7D6",X"00D3D1",X"03D5D4",X"07D9D8",X"01D1D3",X"03CED4",X"11D6DE",X"14D3DD",X"18D0DA",X"25DAE5",X"46B7BB",X"112836",X"000009",X"C7B142",X"F4E74D",X"8C8200",X"060700",X"00000B",X"90727A",X"FCF0FE",X"FBFDFF",X"F6F9FF",X"FFFCFD",X"FFF4F0",X"FFFEFF",X"F8FFFF",X"FFFCFF",X"FDFBFC",X"FFFCCC",X"D8C046",X"E1B924",X"AD881E",X"140200",X"040404",X"512228",X"A22B63",X"B31B70",X"C11577",X"D4077E",X"AC0B6B",X"FFD4FA",X"FCFFFF",X"F7FFFF",X"FFFEFF",X"FFFAFD",X"FFFBFC",X"FEFFFF",X"F8FFFF",X"FCFFFF",X"FFFCFB",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"F3F3F3",X"39363D",X"040001",X"2F2523",X"211000",X"230715",X"240C0A",X"1B080A",X"1E1504",X"26150D",X"2C1817",X"110000",X"ECE0E2",X"FFFCFD",X"FEFFFF",X"FCFFFF",X"F8FAF7",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"F5FFF1",X"FFFAFF",X"FFF8FF",X"C0CEF3",X"0023A2",X"156CBB",X"0D6AC7",X"186DE2",X"0F68E0",X"0966DF",X"0065D2",X"076BDA",X"006BD3",X"1B6ACF",X"004FDE",X"BDD1F4",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FDFDFD",X"F7FFFD",X"8F90BE",X"010200",X"271E15",X"0B0300",X"160F00",X"777300",X"CBC82D",X"F1DD2E",X"E0D018",X"E8D900",X"E5CF00",X"EBDC5B",X"F4FBD1",X"F8FFFD",X"FFF8FF",X"FEFFFF",X"FDFBFC",X"FFFCFE",X"F9F5FF",X"FCFFFF",X"FDFFE4",X"E0E281",X"DCDB45",X"DEC67E",X"83804D",X"080500",X"080000",X"290918",X"260008",X"1E252F",X"48BFAB",X"15D29A",X"0CD090",X"0EC585",X"39C598",X"024D38",X"0D0000",X"9D1E25",X"DD0615",X"D40000",X"ED0707",X"E80809",X"DE0A09",X"E8030A",X"F2000E",X"D50D17",X"98150D",X"1D0002",X"073C28",X"28C192",X"29D7A4",X"098C6A",X"003E23",X"001002",X"0C0001",X"CABE68",X"D9D267",X"CDC771",X"857963",X"110004",X"2F080D",X"2B0009",X"32002A",X"0A0614",X"263C6B",X"3361AF",X"2961B8",X"2165AE",X"2B71A5",X"274C69",X"34313C",X"291023",X"2D0020",X"5A0044",X"85005E",X"BA1782",X"C20D78",X"C6026E",X"C50067",X"C80772",X"C4006B",X"D00379",X"C10F71",X"A42364",X"6C223D",X"260301",X"0E0000",X"430000",X"B86C2E",X"734708",X"030D02",X"170420",X"2B6646",X"0B6F2F",X"146B41",X"065526",X"13743F",X"085727",X"001400",X"060918",X"08000E",X"9C5E47",X"E76F23",X"E06B1C",X"EA6C20",X"E56619",X"DF6C19",X"BB610B",X"894401",X"420A00",X"240000",X"000900",X"120718",X"361F31",X"6D5D4E",X"8F7F5D",X"A18061",X"966D4D",X"92713E",X"907057",X"835E43",X"6C4F3F",X"483A3A",X"0D0001",X"140000",X"040005",X"0F233E",X"040007",X"D6D3E4"),
(X"FFFAFF",X"758D8D",X"008165",X"2DC6AA",X"0FB698",X"14C7A7",X"00BE9F",X"24D4BF",X"27897A",X"000E0E",X"040003",X"432616",X"74471E",X"682400",X"5A0800",X"4C0000",X"540600",X"591A00",X"7C3600",X"C45F0D",X"F17D26",X"F9872F",X"FC8622",X"F57300",X"FE730C",X"FE7C0C",X"F88005",X"F07D00",X"FB830B",X"F67C19",X"EE8534",X"CA782F",X"9A7B5F",X"3B200F",X"0B0000",X"080C0F",X"001114",X"043836",X"0D5853",X"116661",X"0C5D57",X"085A58",X"045357",X"055355",X"115B5C",X"02514E",X"055B5A",X"005B5B",X"105457",X"0F585F",X"0E5D6A",X"035968",X"045A69",X"03565E",X"0E5A5A",X"115A53",X"235B5A",X"1A4649",X"092229",X"050E15",X"02070A",X"000806",X"001009",X"00130C",X"005768",X"04808C",X"26B5BD",X"33D8DC",X"20D9DC",X"0BD5D9",X"05D6DD",X"00CDD7",X"02D9DB",X"09DDE0",X"04D4D8",X"03CED2",X"09D4D8",X"07D5D5",X"07D9D8",X"00D1CF",X"07D9D8",X"08DAD9",X"06D6D8",X"07D2D8",X"0DD2DA",X"0AC9D3",X"0DC5CF",X"17CCD7",X"49BABE",X"1A313F",X"060610",X"A99324",X"F4E74D",X"E6DC58",X"64652B",X"00000B",X"5F4149",X"FDF1FF",X"FAFCFF",X"F7FAFF",X"FFF9FA",X"FFFCF8",X"FCFAFB",X"F4FBFF",X"FFFBFF",X"FFFDFE",X"FFF9C9",X"D0B83E",X"DEB621",X"E9C45A",X"84724C",X"040404",X"35060C",X"830C44",X"BC2479",X"B10567",X"E2158C",X"AC0B6B",X"F6BCE2",X"F6FAFD",X"F4FEFF",X"FFFDFF",X"FFFAFD",X"FFFCFD",X"FEFFFF",X"F8FFFF",X"FCFFFF",X"FFFCFB",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"F3F3F3",X"36333A",X"060203",X"070000",X"110000",X"140006",X"160000",X"0D0000",X"090000",X"0D0000",X"120000",X"0D0000",X"EADEE0",X"FFFEFF",X"F9FAFE",X"F9FDFE",X"FEFFFD",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"F8FFF4",X"FFF9FF",X"FFFBFF",X"CAD8FD",X"0D3AB9",X"237AC9",X"0F6CC9",X"0F64D9",X"0D66DE",X"0865DE",X"046EDB",X"066AD9",X"036ED6",X"2A79DE",X"0156E5",X"B7CBEE",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"F7FFFD",X"9E9FCD",X"000100",X"0B0200",X"766E3D",X"C2BB60",X"DDD951",X"E2DF44",X"E5D122",X"DCCC14",X"E3D400",X"E9D300",X"DECF4E",X"FAFFD7",X"F6FFFB",X"FDF2FF",X"FDFEFF",X"FFFEFF",X"FFFDFF",X"FFFCFF",X"FCFFFF",X"FDFFE4",X"F9FB9A",X"CAC933",X"7F671F",X"0C0900",X"171401",X"261A1E",X"432332",X"410D23",X"00010B",X"229985",X"19D69E",X"00C181",X"0BC282",X"37C396",X"26715C",X"100100",X"8D0E15",X"E30C1B",X"DE0500",X"E50000",X"DC0000",X"DB0706",X"E9040B",X"F1000D",X"D50D17",X"9B1810",X"29090E",X"0B402C",X"21BA8B",X"14C28F",X"40C3A1",X"50B095",X"0B3B2D",X"120107",X"746812",X"A49D32",X"342E00",X"0D0100",X"1B010E",X"4B2429",X"582836",X"3D0A35",X"120E1C",X"000C3B",X"053381",X"2A62B9",X"1559A2",X"003367",X"000825",X"010009",X"240B1E",X"501C43",X"84276E",X"9D1776",X"B91681",X"BB0671",X"C5016D",X"CE0470",X"C2016C",X"D4087B",X"C80071",X"C00E70",X"7F003F",X"400011",X"2B0806",X"2F1D0F",X"A86249",X"CF8345",X"A5793A",X"000A00",X"0B0014",X"023D1D",X"056929",X"085F35",X"075627",X"005E29",X"206F3F",X"062810",X"070A19",X"120318",X"9B5D46",X"ED7529",X"E77223",X"E96B1F",X"EA6B1E",X"E87522",X"E48A34",X"D18C49",X"A56D48",X"764439",X"000600",X"24192A",X"2D1628",X"0D0000",X"5B4B29",X"AE8D6E",X"986F4F",X"866532",X"8D6D54",X"8E694E",X"896C5C",X"9E9090",X"78696C",X"594441",X"272028",X"00112C",X"040007",X"D5D2E3"),
(X"FFFCF9",X"839796",X"008268",X"2BC1A6",X"0EB798",X"08C89F",X"0BCBA4",X"2CBBA7",X"184629",X"000302",X"220B25",X"0E0012",X"150015",X"15000C",X"190012",X"1D0020",X"1B000E",X"0E000E",X"0A0000",X"190400",X"5C3E1C",X"9C6F45",X"C3773B",X"FB8C3B",X"F2720D",X"FC7607",X"FF7A00",X"FD7800",X"FA7902",X"F6790B",X"F98315",X"F98A16",X"FF851E",X"D66B19",X"7F3603",X"1D0000",X"0E0100",X"0D0D0F",X"1D1D25",X"323139",X"1B5758",X"1C605F",X"125E5A",X"05554C",X"0E5E53",X"08554F",X"0D585B",X"095660",X"02625E",X"005F54",X"046552",X"005E48",X"086552",X"015B51",X"0A6061",X"0B5E66",X"034E53",X"0E5C60",X"105B5E",X"094D4C",X"003431",X"001D1F",X"001720",X"001320",X"000704",X"000808",X"071619",X"2A474D",X"559096",X"58BEC0",X"35C6C1",X"23CDC4",X"06C7D0",X"0BCDD7",X"09CFD8",X"0ED8E4",X"09D4E2",X"07D5E3",X"0BD8E9",X"08D7E9",X"0CD5DF",X"08D2DE",X"06D1DF",X"08D3E2",X"06D1E0",X"04CDDD",X"0BD3E3",X"16DEED",X"28BCBE",X"0F343D",X"000200",X"AFA61D",X"F4F52D",X"F8E71E",X"E1CF31",X"7A6F00",X"3F1C08",X"FFF1E7",X"FFFDFF",X"FEF8FF",X"F7F9F8",X"F1FFF6",X"F5FFFD",X"FBFFFF",X"FAFCF1",X"FDFDFF",X"FFFFF1",X"E7D275",X"D6B506",X"E7C406",X"E4CB3B",X"756808",X"150000",X"36130F",X"7D194B",X"C7197B",X"E11171",X"D10662",X"E46CAA",X"FBFFFD",X"F3FBFD",X"FCFEFD",X"FFFFFB",X"FFFFFD",X"FEFFFF",X"FCFFFF",X"FFFFFF",X"FFFDFC",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"F3F3F3",X"38263C",X"6A5A26",X"988121",X"998400",X"988401",X"7C6D00",X"776900",X"5B5000",X"5F4C00",X"6D5A00",X"605005",X"F4EBC4",X"FFFDF4",X"FAFBFD",X"F9FAFF",X"FEFDFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FCFFF1",X"F9F7FA",X"F9FCF5",X"BCD9F9",X"0A44CA",X"187AE5",X"0570E2",X"0169E4",X"0A7EE3",X"006BD8",X"0074DF",X"006EE2",X"0070E0",X"1F76DD",X"0059DE",X"B6D8FD",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFBF4",X"DED9B9",X"7D7812",X"CAC134",X"F0DE4C",X"EEDC22",X"E4D405",X"E8D807",X"EADC07",X"E5CF00",X"DECF1C",X"DED31F",X"DDCF14",X"FAFF93",X"F6FFF2",X"FFFBF8",X"F9FBFA",X"FFFFF5",X"FDFBEE",X"FFFFFB",X"F5F8FF",X"F5F4FC",X"F2E5DF",X"715D44",X"000800",X"2E1116",X"470019",X"A10D57",X"B82365",X"710F36",X"050B0B",X"1E8768",X"27D29D",X"09CA87",X"09CB82",X"20B37D",X"004126",X"0E0000",X"811D1F",X"BA171C",X"D2151B",X"D00A17",X"CB0713",X"CB0D17",X"D10812",X"DA0313",X"C80C1A",X"A00E11",X"2F0007",X"001009",X"37B58F",X"24DCA6",X"0AC78F",X"22CF9A",X"066E4D",X"000400",X"090B08",X"030500",X"250D0D",X"5C114C",X"90046D",X"B70371",X"CB167D",X"A70068",X"6B003F",X"2A0024",X"1D1F34",X"384A54",X"252241",X"1A0036",X"3E003C",X"78094D",X"A50A70",X"BE157A",X"C4076D",X"C30061",X"D0026F",X"CD0478",X"C30279",X"BC0078",X"C31463",X"B41C65",X"90235C",X"5A223B",X"210900",X"2E0700",X"4C0000",X"DA5333",X"E56617",X"F58030",X"C17045",X"0E0004",X"12041D",X"063E1B",X"1A7235",X"1E7042",X"005921",X"0F7438",X"197137",X"1D4925",X"000A03",X"0D0709",X"7E4A32",X"D96C31",X"F16E04",X"FA720F",X"F2670C",X"E75C00",X"FF7012",X"F3630C",X"ED6517",X"ED722C",X"BD5B10",X"661300",X"2D0000",X"110D01",X"303531",X"655558",X"816456",X"957D4D",X"907250",X"A57B51",X"9F7851",X"937B5F",X"9F8D75",X"A58A6D",X"977E60",X"3D311B",X"281C04",X"D0C9B7"),
(X"FFFEFB",X"899D9C",X"03856B",X"28BEA3",X"10B99A",X"02C299",X"18D8B1",X"0E9D89",X"001100",X"000807",X"220B25",X"210825",X"412941",X"38162F",X"3D1436",X"3F1642",X"451A38",X"2C142C",X"130409",X"1A0500",X"190000",X"270000",X"8B3F03",X"E27322",X"F97914",X"FF7B0C",X"FF7A00",X"FF7D00",X"F97801",X"F87B0D",X"F98315",X"EA7B07",X"EF7009",X"F48937",X"D68D5A",X"7D5740",X"0A0000",X"000002",X"0B0B13",X"000007",X"003738",X"0E5251",X"105C58",X"0E5E55",X"07574C",X"125F59",X"0B5659",X"014E58",X"01615D",X"005E53",X"005E4B",X"05644E",X"096653",X"086258",X"075D5E",X"075A62",X"125D62",X"126064",X"0E595C",X"135756",X"1F5653",X"234C4E",X"1D3F48",X"0B2B38",X"000F0C",X"000A0A",X"011013",X"00080E",X"00141A",X"006365",X"1BACA7",X"23CDC4",X"1EDFE8",X"10D2DC",X"04CAD3",X"08D2DE",X"00C9D7",X"01CFDD",X"02CFE0",X"00CFE1",X"0ED7E1",X"05CFDB",X"04CFDD",X"06D1E0",X"00CAD9",X"00C4D4",X"04CCDC",X"0ED6E5",X"21B5B7",X"092E37",X"000200",X"B7AE25",X"F2F32B",X"D8C700",X"F9E749",X"D0C551",X"5F3C28",X"C8B6AC",X"FFFAFE",X"FFFCFF",X"FDFFFE",X"EEFEF3",X"F5FFFD",X"F9FEFF",X"FFFFF6",X"FCFCFF",X"FEF8EA",X"F7E285",X"DDBC0D",X"D4B100",X"E7CE3E",X"C5B858",X"270907",X"1D0000",X"61002F",X"B80A6C",X"F12181",X"C9005A",X"EE76B4",X"EBF1ED",X"F6FEFF",X"FDFFFE",X"FFFFFB",X"FFFFFD",X"FEFFFF",X"FCFFFF",X"FFFFFF",X"FFFDFC",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"F3F3F3",X"110015",X"948450",X"F0D979",X"E1CC3D",X"E4D04D",X"D1C245",X"E0D267",X"C2B74B",X"CDBA54",X"DFCC6D",X"C1B166",X"FFFCD5",X"FFFEF5",X"FEFFFF",X"FEFFFF",X"FEFDFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FCFFF1",X"FBF9FC",X"FEFFFA",X"BAD7F7",X"0C46CC",X"1274DF",X"0570E2",X"0870EB",X"077BE0",X"006FDC",X"017AE5",X"0978EC",X"0173E3",X"166DD4",X"0053D8",X"ACCEF3",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFF8",X"FDF8D8",X"E6E17B",X"E1D84B",X"DAC836",X"E0CE14",X"E4D405",X"E1D100",X"ECDE09",X"E5CF00",X"DDCE1B",X"DCD11D",X"DDCF14",X"E2EA7B",X"F4FFF0",X"FFFBF8",X"F9FBFA",X"FFFFF6",X"FFFEF1",X"FFFFFB",X"FCFFFF",X"FFFEFF",X"FFF5EF",X"5E4A31",X"000900",X"492C31",X"7D1C4F",X"B6226C",X"AF1A5C",X"8D2B52",X"000202",X"147D5E",X"26D19C",X"04C582",X"03C57C",X"2EC18B",X"004328",X"0B0000",X"791517",X"B8151A",X"C5080E",X"CE0815",X"D30F1B",X"CD0F19",X"D00711",X"E10A1A",X"D41826",X"AA181B",X"440E1C",X"000700",X"189670",X"28E0AA",X"03C088",X"1ECB96",X"369E7D",X"000B05",X"1F211E",X"282A15",X"351D1D",X"6A1F5A",X"AD218A",X"BF0B79",X"BD086F",X"B70D78",X"89135D",X"40073A",X"06081D",X"000D17",X"00001B",X"290545",X"661864",X"922367",X"AD1278",X"BF167B",X"C5086E",X"CB0069",X"CB006A",X"C60071",X"C5047B",X"C2047E",X"BD0E5D",X"A9115A",X"670033",X"2A000B",X"120000",X"77502F",X"C56B46",X"E76040",X"DF6011",X"F88333",X"C57449",X"0A0000",X"0A0015",X"0C4421",X"11692C",X"1D6F41",X"076028",X"1A7F43",X"096127",X"295531",X"112019",X"040000",X"4A1600",X"CE6126",X"E96600",X"EB6300",X"F66B10",X"F56A0D",X"F8690B",X"E75700",X"ED6517",X"EE732D",X"E7853A",X"BE6B41",X"5B2D1D",X"0A0600",X"404541",X"28181B",X"634638",X"7C6434",X"7E603E",X"9B7147",X"956E47",X"897155",X"99876F",X"9E8366",X"A68D6F",X"736751",X"756951",X"EAE3D1"),
(X"FEFFFA",X"779A93",X"039878",X"15C0A0",X"07C19C",X"0CCA9E",X"34C5A6",X"2C605E",X"000600",X"2A042B",X"61045F",X"830F8C",X"91139B",X"900B98",X"9B18A6",X"850C99",X"94088D",X"82058D",X"6E047E",X"4C0054",X"34003E",X"190021",X"130000",X"482B0B",X"B76E39",X"E7873D",X"FC7C1B",X"FF7308",X"FE7107",X"F77307",X"FF7E0B",X"FF7A00",X"FF8211",X"EF7102",X"FC8414",X"F58A20",X"C66E15",X"541700",X"200000",X"150000",X"1A0600",X"0A0600",X"102423",X"29565C",X"1C5860",X"10575B",X"055556",X"0B605D",X"005D5A",X"005A5A",X"035A61",X"0B5D68",X"0C5B68",X"085863",X"03585F",X"045B62",X"06535D",X"065D64",X"005F5F",X"006059",X"005D53",X"0C5953",X"195659",X"174B56",X"00433A",X"002F29",X"00201E",X"001518",X"000E14",X"00050B",X"000C13",X"2C4349",X"5195A2",X"51A8B1",X"4AC0C2",X"39CECC",X"16C3BD",X"14CDC8",X"10CCCB",X"0ECACB",X"01D3D2",X"00CECF",X"00D1D4",X"03D6DD",X"02D3DA",X"00CFD9",X"08D4DD",X"10DAE4",X"30B5BA",X"152535",X"0D0200",X"938626",X"F1F362",X"FEE854",X"FAE25E",X"E1D461",X"989163",X"919475",X"FEFFFA",X"FFFAFF",X"FFF9FD",X"FEFFFD",X"F9FEF8",X"FEFDFB",X"FCFCFC",X"FCFFFF",X"FAFCF1",X"EBDFA5",X"DAB934",X"EABE03",X"E6BF02",X"E1C120",X"BD9B3A",X"000600",X"0D0E10",X"380B10",X"972D5B",X"AF075F",X"D13888",X"FFD0FF",X"FFFEFF",X"FCFFFD",X"F8FFF9",X"F7FFF9",X"FEFFFF",X"FFFDFF",X"FFFDFF",X"FFFDFE",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"F3F3F3",X"101221",X"908D18",X"E8CA36",X"E8C104",X"E4BA06",X"EDC01C",X"F3BF1E",X"F2B715",X"E4C709",X"E8D111",X"CCBD22",X"FFF6AB",X"FCFAEB",X"F8FCFD",X"F7F8FC",X"FFFCFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFC",X"FBFAF8",X"F8FFF4",X"B8DEF5",X"0E50C1",X"0F71DC",X"006DCF",X"0170C9",X"0065C5",X"006DD6",X"036BDA",X"0B66D9",X"0C64CE",X"296EC9",X"165BC0",X"AECDEA",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"F7F6FF",X"FFFFD2",X"D4D062",X"D4CF04",X"EEDC22",X"E4D109",X"EED910",X"E3D101",X"E1D505",X"F4D900",X"E3D512",X"E8D821",X"F5CE04",X"ECD956",X"FEFFEB",X"FFF4FE",X"FEFEFF",X"FFFFFF",X"FFFFFA",X"FBFEF7",X"F5F9FA",X"FDF9FF",X"FCECFF",X"876C8F",X"800039",X"C51E7A",X"CC0C7D",X"D2057B",X"C61570",X"6A153F",X"000704",X"1D6D52",X"33CBA2",X"0BCF8F",X"00CD83",X"29D297",X"248164",X"000A02",X"3C201C",X"642B24",X"551A1C",X"5D1C22",X"642329",X"5C2221",X"551E17",X"5F261D",X"632A23",X"5B2421",X"250510",X"122B25",X"239574",X"1DD29D",X"00CC8D",X"04D996",X"36C897",X"275342",X"040011",X"132227",X"2D1F2C",X"972C64",X"B90664",X"CA0D74",X"BB076A",X"CB1172",X"C9176F",X"90105D",X"500033",X"4A001F",X"6C002E",X"9F0A5C",X"BF0776",X"CF0278",X"B1006A",X"BC0466",X"CE0B6B",X"D30A70",X"C0006D",X"B60C6F",X"B4226B",X"A9295C",X"911E45",X"41081B",X"040000",X"3D3119",X"8A421C",X"DD6028",X"FB7221",X"E36801",X"F36F0B",X"DE762F",X"B77360",X"040006",X"000A05",X"014D1C",X"095F22",X"045D2F",X"136A35",X"00622B",X"126B35",X"30673D",X"415E48",X"000902",X"190000",X"AC5D4E",X"D67C3E",X"D87534",X"E56420",X"F45406",X"FF6504",X"FA7204",X"EF6B00",X"F96505",X"E36000",X"FC6D1E",X"F17339",X"9A5220",X"150000",X"31281F",X"080000",X"5A4F4B",X"846A5D",X"A77E62",X"7C4E2A",X"866242",X"927356",X"9C7652",X"AE8157",X"A27349",X"76623F",X"EBDCBB"),
(X"FEFFFA",X"8EB1AA",X"0EA383",X"11BC9C",X"02BC97",X"0FCDA1",X"2ABB9C",X"002E2C",X"000500",X"2B052C",X"761974",X"8C1895",X"83058D",X"8A0592",X"8B0896",X"7E0592",X"94088D",X"8C0F97",X"801690",X"77227F",X"481152",X"200528",X"210C0B",X"190000",X"681F00",X"D07026",X"FF8726",X"FE6D02",X"FC6F05",X"F77307",X"FC7603",X"FF7700",X"F67807",X"F97B0C",X"ED7505",X"F68B21",X"E99138",X"CD9051",X"7F5839",X"371C15",X"110000",X"040000",X"000E0D",X"001C22",X"003941",X"0B5256",X"136364",X"0C615E",X"00615E",X"005A5A",X"055C63",X"035560",X"0F5E6B",X"085863",X"095E65",X"035A61",X"105D67",X"0E656C",X"016565",X"00645D",X"015E54",X"095650",X"165356",X"164A55",X"1C5F56",X"154E48",X"1D4745",X"173336",X"04171D",X"000F15",X"000D14",X"00080E",X"001724",X"004E57",X"178D8F",X"17ACAA",X"0DBAB4",X"1AD3CE",X"1BD7D6",X"18D4D5",X"01D3D2",X"00D2D3",X"00D1D4",X"00D0D7",X"00CFD6",X"00CDD7",X"05D1DA",X"0ED8E2",X"29AEB3",X"0D1D2D",X"0A0000",X"908323",X"EEF05F",X"DFC935",X"BCA420",X"ADA02D",X"5E5729",X"8E9172",X"FEFFFA",X"FAF3FA",X"FFF9FD",X"FEFFFD",X"F6FBF5",X"FFFFFD",X"FBFBFB",X"F8FCFF",X"FFFFF6",X"FEF2B8",X"DBBA35",X"E9BD02",X"E0B900",X"E7C726",X"E7C564",X"7D8465",X"000002",X"33060B",X"5E0022",X"C82078",X"AA1161",X"ECA4D6",X"FEFCFF",X"FBFFFC",X"F8FFF9",X"F7FFF9",X"FEFFFF",X"FFFDFF",X"FFFDFF",X"FFFDFE",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"F3F3F3",X"181A29",X"7F7C07",X"E9CB37",X"E9C205",X"ECC20E",X"F1C420",X"F0BC1B",X"F4B917",X"D9BC00",X"D9C202",X"C6B71C",X"FFF6AB",X"FFFFF1",X"FCFFFF",X"FCFDFF",X"FFFDFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FCFBF9",X"F9F8F6",X"F7FFF3",X"B5DBF2",X"1153C4",X"1577E2",X"0171D3",X"0473CC",X"0071D1",X"0774DD",X"036BDA",X"146FE2",X"166ED8",X"2E73CE",X"0F54B9",X"B3D2EF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"F8F7FF",X"FFFFD6",X"F1ED7F",X"D2CD02",X"E0CE14",X"F5E21A",X"DFCA01",X"E5D303",X"DBCF00",X"FDE200",X"E3D512",X"E7D720",X"EFC800",X"EBD855",X"FAFCE7",X"FFF4FE",X"FBFBFF",X"F8F8FA",X"FEFFF9",X"FEFFFA",X"FCFFFF",X"FFFCFF",X"FFF7FF",X"D8BDE0",X"94094D",X"C31C78",X"C30374",X"D2057B",X"BC0B66",X"69143E",X"000E0B",X"0C5C41",X"1CB48B",X"0ED292",X"00C77D",X"1AC388",X"137053",X"000901",X"2C100C",X"3B0200",X"350000",X"350000",X"350000",X"2E0000",X"2B0000",X"2C0000",X"2B0000",X"300000",X"150000",X"00120C",X"178968",X"19CE99",X"00CA8B",X"06DB98",X"30C291",X"1D4938",X"030010",X"031217",X"080007",X"841951",X"C61371",X"BA0064",X"C41073",X"B90060",X"B9075F",X"A32370",X"752258",X"732348",X"902052",X"AD186A",X"BE0675",X"D1047A",X"C2117B",X"BA0264",X"C90666",X"CA0167",X"C70774",X"C1177A",X"A8165F",X"860639",X"5E0012",X"3F0619",X"050000",X"6B5F47",X"D8906A",X"E76A32",X"F46B1A",X"EB7009",X"FC7814",X"D46C25",X"6C2815",X"060108",X"07221D",X"0B5726",X"12682B",X"076032",X"237A45",X"046730",X"07602A",X"1C5329",X"27442E",X"000700",X"30120A",X"A05142",X"AD5315",X"B14E0D",X"E86723",X"FF6618",X"FF6504",X"F76F01",X"EC6800",X"FC6808",X"F47105",X"F16213",X"E96B31",X"C47C4A",X"8C7452",X"070000",X"120608",X"1F1410",X"795F52",X"AA8165",X"9F714D",X"B38F6F",X"A7886B",X"6B4521",X"92653B",X"AE7F55",X"6A5633",X"DBCCAB"),
(X"F8FBF4",X"90CEBF",X"05AA88",X"14BBA1",X"06B596",X"26BD9E",X"348274",X"010007",X"1D0D34",X"480353",X"820784",X"920298",X"A00BA5",X"980498",X"860085",X"941998",X"A51CAA",X"880099",X"8C009A",X"9B0D9D",X"951495",X"6E0878",X"3F0048",X"34002E",X"080004",X"623E26",X"D58747",X"F2771A",X"FF7307",X"FF7A0A",X"FC7404",X"FC6E02",X"FD7708",X"F97200",X"FF7802",X"FF7A00",X"FE8007",X"FB871A",X"F78E33",X"CD6C1F",X"8B3A0B",X"561400",X"290000",X"110000",X"14100D",X"09160F",X"0C281C",X"294F40",X"17515C",X"125158",X"115554",X"09544D",X"0C5D54",X"085F56",X"09625C",X"045F5A",X"005556",X"055F60",X"046262",X"06655F",X"045F56",X"015B51",X"08615B",X"096562",X"014A5D",X"0A5966",X"085D64",X"085E5F",X"085452",X"003838",X"001F20",X"001416",X"000907",X"000305",X"000107",X"00000B",X"172532",X"395B65",X"51888D",X"62A8AA",X"43BDCC",X"47C6D5",X"3EC6D4",X"30C4D2",X"25C6D0",X"19C6CD",X"13C9CD",X"19D2D5",X"3FBAB5",X"0F313B",X"000707",X"565541",X"706851",X"2D0F05",X"140000",X"0B0000",X"240000",X"6D4649",X"EFE0E7",X"FAFDFF",X"FEFFFF",X"FFFAFC",X"FFF8FB",X"FFFCFF",X"FFFFF6",X"F6F8F7",X"F9FBFF",X"FFFDF2",X"DFC76F",X"DFB513",X"EABF1A",X"E9C648",X"D3B847",X"6F8959",X"0A001A",X"1C001A",X"000200",X"702858",X"AA0262",X"FF8BCD",X"FFEFFB",X"FFF9FB",X"F9FFFA",X"F8FFFA",X"FEFEFE",X"FFFCFF",X"FFFDFF",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"F3F3F3",X"1C203B",X"7A7800",X"F8D63F",X"E9C109",X"E3C40A",X"D5BE0E",X"DBC300",X"E1BE00",X"EDB915",X"E7C00B",X"D0B726",X"FFF1B8",X"FFFAFF",X"FCFFFF",X"FCFFF8",X"FFFCF9",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFCFF",X"FFFDFF",X"F9FFFF",X"BCD5FD",X"1F4BAE",X"336FE1",X"2466D6",X"296DD0",X"3271BE",X"2B62B4",X"3160AE",X"446BB0",X"395E92",X"3C597B",X"061E40",X"B9C0C8",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"F9FFFF",X"FAF9E7",X"F4EAAF",X"D0CB0D",X"ECDF04",X"E6D30B",X"F1E20D",X"DDD100",X"E2D400",X"EDDA00",X"E1D409",X"DECA13",X"E9C70D",X"E2D531",X"E6F49F",X"F6FFF5",X"FFFEFF",X"FCFBFF",X"FCFCFF",X"FCFFFF",X"FCFFFB",X"FEFDF8",X"FFF6F7",X"E9D8E2",X"960852",X"CD1B7B",X"BC006D",X"CA0076",X"D70D79",X"A0175F",X"1E000F",X"1E222B",X"3CB69F",X"28CFA3",X"02C488",X"22C896",X"006E51",X"001C0F",X"001608",X"000F02",X"000F0B",X"001A11",X"002315",X"001E0E",X"001F0E",X"001E0C",X"001E0C",X"003420",X"00442B",X"003C1C",X"03A171",X"21DCA5",X"00C489",X"03D190",X"25C690",X"0B573B",X"00070D",X"13031E",X"280324",X"2F0013",X"7D2243",X"BC206A",X"CD0A73",X"C70170",X"C10F65",X"D11B89",X"C3067E",X"C6026E",X"CA0668",X"C80A6E",X"BC066B",X"B90568",X"C80480",X"C90077",X"DD1180",X"C80968",X"B21861",X"781848",X"310E26",X"10141D",X"0D2B23",X"000807",X"00080B",X"403635",X"7D5347",X"B46F52",X"CD7649",X"DB7B48",X"BD7948",X"7A583C",X"0A0000",X"000F04",X"03471E",X"075F22",X"105F28",X"076334",X"055928",X"0E6C3A",X"095F32",X"1E5737",X"0D3221",X"00070D",X"23102E",X"470D3D",X"1B0008",X"140000",X"835F45",X"CC8454",X"DE6828",X"F15F12",X"F36209",X"E35D00",X"F9711D",X"EC5703",X"FF7518",X"F36F0B",X"E6741E",X"973F0F",X"2A0200",X"00020C",X"4D3D3E",X"8E756E",X"B69785",X"AF8B71",X"9E7557",X"855735",X"906240",X"8C6141",X"927F61",X"F4E6CB"),
(X"FEFFFA",X"80BEAF",X"03A886",X"1BC2A8",X"0AB99A",X"27BE9F",X"004D3F",X"020008",X"110128",X"5A1565",X"931895",X"89008F",X"9B06A0",X"990599",X"920891",X"8D1291",X"99109E",X"9105A2",X"9202A0",X"900292",X"860586",X"811B8B",X"6A2173",X"390033",X"140710",X"1C0000",X"AA5C1C",X"F2771A",X"FD7004",X"FE7606",X"FC7404",X"FF7509",X"F87203",X"FE7704",X"FC7400",X"FF7C01",X"F77900",X"EE7A0D",X"EB8227",X"DD7C2F",X"D28152",X"C2805D",X"6D402D",X"140000",X"030000",X"08150E",X"001105",X"002617",X"07414C",X"14535A",X"115554",X"135E57",X"004E45",X"045B52",X"015A54",X"09645F",X"045A5B",X"045E5F",X"005E5E",X"04635D",X"045F56",X"005A50",X"055E58",X"05615E",X"0D5669",X"0B5A67",X"01565D",X"065C5D",X"0F5B59",X"195555",X"255152",X"1E4042",X"0E2220",X"030E10",X"060B11",X"00010C",X"000613",X"000913",X"001318",X"003C3E",X"00707F",X"0D8C9B",X"1AA2B0",X"1EB2C0",X"25C6D0",X"21CED5",X"1CD2D6",X"25DEE1",X"4CC7C2",X"1B3D47",X"000808",X"050400",X"080000",X"1F0100",X"341817",X"2E1F22",X"5C2926",X"260002",X"D7C8CF",X"FCFFFF",X"F6F7F9",X"FFFBFD",X"FFFAFD",X"FFFAFD",X"FAFCF1",X"FEFFFF",X"FBFDFF",X"FEFAEF",X"E5CD75",X"DDB311",X"F7CC27",X"DDBA3C",X"856A00",X"000D00",X"160726",X"250423",X"020806",X"3B0023",X"A4005C",X"C0387A",X"FEE8F4",X"FDF7F9",X"F9FFFA",X"F8FFFA",X"FEFEFE",X"FFFAFF",X"FFFCFF",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"F3F3F3",X"242843",X"737100",X"E3C12A",X"F4CC14",X"E3C40A",X"E0C919",X"DFC703",X"EBC800",X"F0BC18",X"E2BB06",X"CAB120",X"FFF4BB",X"FFFCFF",X"FAFDFF",X"FBFEF7",X"FFFEFB",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEF7FE",X"FFFDFF",X"F9FFFF",X"B9D2FA",X"1440A3",X"2561D3",X"1355C5",X"1A5EC1",X"104F9C",X"033A8C",X"073684",X"052C71",X"001B4F",X"133052",X"000325",X"BDC4CC",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"F9FFFF",X"FBFAE8",X"FFFABF",X"E3DE20",X"E5D800",X"E9D60E",X"EADB06",X"EDE100",X"F1E306",X"E3D000",X"EDE015",X"E3CF18",X"FFE026",X"E0D32F",X"DCEA95",X"F9FFF8",X"FEFCFF",X"FFFEFF",X"FEFEFF",X"FCFFFF",X"F6FBF5",X"FFFEF9",X"FFFCFD",X"F6E5EF",X"D44690",X"BB0969",X"D11182",X"CB0177",X"CE0470",X"A41B63",X"330824",X"0B0F18",X"2DA790",X"22C99D",X"03C589",X"15BB89",X"38AB8E",X"2A7669",X"3C7668",X"477568",X"48716D",X"4E8D84",X"4B9D8F",X"408E7E",X"4B8B7A",X"508D7B",X"4A8D7B",X"5AA591",X"52A289",X"3CA989",X"22C090",X"13CE97",X"0CD297",X"03D190",X"21C28C",X"2D795D",X"000309",X"352540",X"1F001B",X"240008",X"690E2F",X"BE226C",X"C20068",X"CE0877",X"C6146A",X"CD1785",X"C0037B",X"C90571",X"C60264",X"C00266",X"BD076C",X"C00C6F",X"C3007B",X"CA0078",X"E31786",X"BF005F",X"A0064F",X"530023",X"16000B",X"20242D",X"335149",X"223C3B",X"000508",X"100605",X"240000",X"581300",X"963F12",X"A0400D",X"7D3908",X"1B0000",X"190B08",X"0C261B",X"1D6138",X"146C2F",X"095821",X"015D2E",X"0E6231",X"0F6D3B",X"247A4D",X"1C5535",X"153A29",X"000A10",X"190624",X"3B0131",X"2C0719",X"250908",X"5A361C",X"762E00",X"E06A2A",X"FF7225",X"EB5A01",X"FC7617",X"E9610D",X"FD6814",X"EE5B00",X"F97511",X"CF5D07",X"CF7747",X"572F25",X"00020C",X"100001",X"523932",X"A38472",X"B59177",X"865D3F",X"B18361",X"875937",X"966B4B",X"6E5B3D",X"E6D8BD"),
(X"FFFEFD",X"7BC9B9",X"05AE8D",X"28B5A5",X"2CB5A3",X"369086",X"00070B",X"0B0811",X"5A0058",X"9E1891",X"99008C",X"930190",X"910896",X"92018E",X"97008A",X"9A028B",X"A00191",X"950095",X"900199",X"8D038E",X"92048C",X"960996",X"860C92",X"731180",X"1C002E",X"0C000B",X"432405",X"CF8031",X"FA8211",X"FA7900",X"F87800",X"FB7408",X"FD7700",X"F97400",X"FC7A0C",X"F6770C",X"FA7C0D",X"FC7905",X"FF7A02",X"FD7100",X"FF7508",X"F6760B",X"F98927",X"D47521",X"742800",X"290000",X"160000",X"130212",X"0F0800",X"0C1002",X"183023",X"245248",X"1B5850",X"10574F",X"145F58",X"0F5C54",X"005B55",X"05615E",X"025A5B",X"07565A",X"105C5C",X"075756",X"005454",X"0A6E6E",X"035C58",X"065C59",X"085C5C",X"085859",X"0C5A5C",X"035153",X"0D5B5D",X"0C5A5C",X"125B52",X"054C44",X"003B34",X"002F2D",X"00292A",X"002026",X"00111A",X"000712",X"020808",X"000302",X"000404",X"102526",X"264643",X"3D6662",X"406F67",X"4C7F76",X"608D93",X"252233",X"040004",X"660C3F",X"A31464",X"AF0369",X"B8117A",X"BB147D",X"C41270",X"AA0259",X"FFA1DB",X"FFEDFF",X"EDFFFD",X"FBFFFD",X"FBF2F7",X"FFFEFF",X"FFFCFF",X"FFFCF9",X"FCFFFF",X"FAFFFC",X"F6ECBB",X"E5C860",X"D0B94F",X"544F0B",X"02000E",X"00071F",X"10427F",X"225CAE",X"001D56",X"01011B",X"4A061F",X"891333",X"F1CEE2",X"FFF9FF",X"FEFFFA",X"F9FEF8",X"FFFFFD",X"FFFAFF",X"FFFDFF",X"FBFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FEFEFE",X"FEFEFE",X"FFFFFF",X"F4F4F4",X"241654",X"786700",X"F0C238",X"EEBF00",X"E6C500",X"DDC606",X"DEC400",X"E6C300",X"F4C311",X"DEB900",X"C6AF13",X"FCEEAD",X"FFFEFD",X"FCFFFF",X"FAFDF6",X"FFFEFB",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFDFF",X"F9F4F8",X"FEFEFF",X"C7CDD9",X"000400",X"202D35",X"020F15",X"010C0E",X"000400",X"000200",X"0C0700",X"070300",X"0A0400",X"090600",X"130300",X"CFC2AF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFDFF",X"FFF1FF",X"FFF7FA",X"F3DB6D",X"E4D403",X"F1D91D",X"EDD80B",X"ECD910",X"E8D41B",X"D7D822",X"E0E33A",X"E1DB61",X"A59C61",X"A48E77",X"7E685B",X"EFF4F0",X"FFFFEF",X"FCFBF6",X"FCFFFF",X"FBFFFF",X"FEFFFD",X"FFFFFA",X"FFFBF9",X"FFF7FD",X"E590BA",X"A60855",X"DA1378",X"D1036F",X"D90A72",X"AA0F5B",X"31001D",X"000507",X"1EAF88",X"13C68F",X"09D492",X"00C282",X"0EC58C",X"1CD19C",X"16C793",X"1CC493",X"1ED39C",X"07BC89",X"26D7A9",X"15C999",X"09C48D",X"15D69D",X"12CF99",X"13C798",X"14D89A",X"0ED094",X"05D091",X"01C88D",X"09D495",X"06D795",X"1CBD87",X"014B30",X"000002",X"4F225B",X"733A89",X"0E0021",X"07000C",X"5F1E49",X"B3237B",X"C30573",X"BD036E",X"C3006D",X"CA0066",X"CC0562",X"C90269",X"D1077F",X"CC0174",X"CC0464",X"CE0070",X"C81974",X"991F5C",X"631B41",X"1C0015",X"000005",X"000D00",X"154422",X"2A703C",X"18633A",X"004529",X"043023",X"000908",X"060000",X"080500",X"000400",X"000500",X"062A1C",X"0A3325",X"124121",X"166E32",X"11652A",X"08521F",X"126F36",X"005D22",X"05672E",X"16693F",X"164A34",X"000E0F",X"020018",X"45185D",X"6C1F87",X"5A1767",X"4C064F",X"3F1140",X"10000B",X"633D2A",X"CB663C",X"EC631D",X"F57011",X"F7630D",X"F9650F",X"EB5E04",X"F56B08",X"FF6E0B",X"F26513",X"BC5B28",X"2D0000",X"261607",X"2F2820",X"5A564D",X"99856D",X"AD865F",X"8A6036",X"896E50",X"9B8E7B",X"150505",X"DBD1D2"),
(X"FAF6F5",X"82D0C0",X"07B08F",X"29B6A6",X"30B9A7",X"116B61",X"00070B",X"120F18",X"861D84",X"900A83",X"99008C",X"9C0A99",X"8D0492",X"960592",X"A10894",X"970088",X"9A008B",X"950095",X"93049C",X"900691",X"90028A",X"910491",X"860C92",X"791786",X"3D1D4F",X"0D000C",X"200100",X"A35405",X"FA8211",X"FF8301",X"FD7D00",X"FD760A",X"FD7700",X"F97400",X"FD7B0D",X"F7780D",X"F97B0C",X"FA7703",X"FF7A02",X"FF7400",X"FE7407",X"F6760B",X"F0801E",X"E38430",X"CD8143",X"AE7957",X"644540",X"0C000B",X"070000",X"000400",X"000900",X"00170D",X"003028",X"00443C",X"034E47",X"17645C",X"04635D",X"005754",X"075F60",X"004E52",X"0B5757",X"095958",X"086262",X"0A6E6E",X"035C58",X"065C59",X"075B5B",X"0D5D5E",X"0F5D5F",X"075557",X"085658",X"045254",X"0E574E",X"0E554D",X"145750",X"1E5A58",X"235657",X"1D464C",X"10313A",X"08232E",X"0B1111",X"020B0A",X"000606",X"00090A",X"000A07",X"00120E",X"000F07",X"00130A",X"000F15",X"070415",X"0F080F",X"6D1346",X"B62777",X"C91D83",X"C21B84",X"BC157E",X"D2207E",X"BA1269",X"CC5F99",X"FFE9FB",X"EBFFFB",X"FBFFFD",X"FFFCFF",X"FCFBFF",X"FCF9FF",X"FFFDFA",X"F9FDFC",X"FBFFFD",X"FEF4C3",X"C7AA42",X"735C00",X"0C0700",X"00000C",X"2C445C",X"3466A3",X"3872C4",X"134079",X"000017",X"4C0821",X"6D0017",X"C5A2B6",X"FFF2FA",X"FFFFFB",X"F8FDF7",X"FDFCFA",X"FFFBFF",X"FFFEFF",X"F7FDFB",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FEFEFE",X"FEFEFE",X"FFFFFF",X"F4F4F4",X"261856",X"786700",X"ECBE34",X"E9BA00",X"DFBE00",X"DAC303",X"E2C800",X"E2BF00",X"DCAB00",X"E4BF00",X"DDC62A",X"FFFBBA",X"FFFBFA",X"FCFFFF",X"F7FAF3",X"FDF9F6",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFCFF",X"FCF7FB",X"FEFEFF",X"C4CAD6",X"000703",X"00060E",X"00060C",X"0D181A",X"141B13",X"434538",X"36311B",X"7D7953",X"A6A06C",X"99965F",X"BAAA76",X"F4E7D4",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFF4FF",X"FFF1F4",X"FBE375",X"DACA00",X"E7CF13",X"DCC700",X"EFDC13",X"FBE72E",X"DCDD27",X"BCBF16",X"666000",X"150C00",X"120000",X"150000",X"DCE1DD",X"FFFAEA",X"F7F6F1",X"FCFFFF",X"FBFFFF",X"FDFFFC",X"FBFAF5",X"FFF9F7",X"FFFBFF",X"FFACD6",X"B0125F",X"D40D72",X"D1036F",X"D1026A",X"B11662",X"32001E",X"000608",X"13A47D",X"16C992",X"00C886",X"0BCF8F",X"0DC48B",X"1CD19C",X"13C490",X"23CB9A",X"0ABF88",X"15CA97",X"13C496",X"19CD9D",X"0CC790",X"03C48B",X"0AC791",X"0EC293",X"12D698",X"09CB8F",X"01CC8D",X"00C68B",X"04CF90",X"07D896",X"24C58F",X"0B553A",X"030305",X"53265F",X"733A89",X"200633",X"07000C",X"43022D",X"A3136B",X"C30573",X"CD137E",X"C90573",X"C90065",X"CC0562",X"CB046B",X"C30071",X"C80070",X"D40C6C",X"DA0A7C",X"B40560",X"8A104D",X"350013",X"12000B",X"1B1E23",X"234230",X"1A4927",X"135925",X"0F5A31",X"0D5236",X"103C2F",X"242E2D",X"0D0503",X"0B0801",X"070F04",X"051000",X"284C3E",X"2C5547",X"2C5B3B",X"0D6529",X"065A1F",X"1C6633",X"0C6930",X"016328",X"096B32",X"196C42",X"073B25",X"00090A",X"010017",X"53266B",X"73268E",X"5F1C6C",X"631D66",X"390B3A",X"22121D",X"1D0000",X"831E00",X"F46B25",X"F87314",X"F5610B",X"FB6711",X"EB5E04",X"EF6502",X"FE6C09",X"EA5D0B",X"E2814E",X"7F4D32",X"100000",X"060000",X"524E45",X"7B674F",X"9F7851",X"A0764C",X"7F6446",X"574A37",X"0E0000",X"DAD0D1"),
(X"FFFDFE",X"7FCCBC",X"00A983",X"25B7A0",X"41B0A0",X"0C2D32",X"11000F",X"2E1E2B",X"6D3272",X"712168",X"812675",X"712273",X"6C1B77",X"7F1581",X"930D8A",X"98088C",X"8F0187",X"920096",X"92019A",X"8F0590",X"930087",X"9C008F",X"9B0096",X"920893",X"801573",X"2A0034",X"0A0004",X"6B360E",X"EA8028",X"FC7F07",X"FB7B00",X"FF7B0C",X"F2780B",X"F47409",X"FF790E",X"FF7605",X"FF7800",X"F87600",X"F77F04",X"F17F05",X"F78008",X"FB830B",X"FB7E06",X"F77500",X"FE7807",X"FF8620",X"EC7A24",X"C0580F",X"933500",X"701E00",X"4A0B00",X"250000",X"0D0000",X"140F16",X"191E22",X"283032",X"1E4847",X"1B4B4F",X"1B5257",X"246166",X"185C5F",X"0D565C",X"01545A",X"015B64",X"03625E",X"06605E",X"035759",X"0B5C5F",X"0B5C5F",X"055E5C",X"01625B",X"006259",X"086061",X"075D5E",X"085C5C",X"0C615E",X"0F615F",X"0A5C58",X"075955",X"095B55",X"0D4F4E",X"0F4C4D",X"0C4348",X"02313B",X"001E2A",X"001A29",X"000C1A",X"000917",X"000907",X"000308",X"030600",X"770342",X"D81274",X"EC027B",X"E5017A",X"EB037D",X"E20892",X"E1017E",X"E22F8A",X"FFD0F8",X"FFFCFF",X"F3FCF9",X"FEFFFF",X"FBFFFF",X"FFFCFF",X"FFFEF6",X"FEFFED",X"F1FCF8",X"F6F4F5",X"A9978D",X"000002",X"042946",X"0043AD",X"0878DC",X"077AD5",X"106AD8",X"1664E2",X"043488",X"08192D",X"000402",X"8B6F86",X"FFEFFD",X"FAF4F6",X"FFFFFB",X"FFFEFF",X"F9F7FA",X"FDFDFF",X"FCFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FEFEFE",X"FEFEFE",X"FFFFFF",X"F4F4F4",X"23262F",X"706C00",X"E1C442",X"E4C014",X"DAB90C",X"DBBA15",X"E8C426",X"E0B318",X"D8B31A",X"CFB311",X"C8B733",X"F9F1B0",X"FEFEF2",X"F9FDFC",X"FFFFFD",X"FFFDFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFDFF",X"FFFFF8",X"FFFEFB",X"E1DBA9",X"817D00",X"A09300",X"CCBD18",X"DACD26",X"C8C311",X"DDD31A",X"E0D116",X"EEE71D",X"EAE118",X"E7E52E",X"EED823",X"FAF79A",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"F5F9EB",X"FFFBFA",X"FFFCF3",X"FFF1C0",X"D6D23B",X"E4DD4F",X"EEE661",X"D3C564",X"B09965",X"6E744E",X"0C0902",X"090100",X"0A0905",X"571942",X"780143",X"F08CAE",X"FFF9FF",X"FFFBFF",X"FCFDFF",X"F7FBFE",X"F9FBF8",X"FFFEFF",X"FFFDFF",X"FFFAFF",X"F7DEF4",X"AF3872",X"CC0E66",X"CE0666",X"C90E67",X"AB1A5B",X"44041E",X"030500",X"2B8965",X"4DC095",X"44C897",X"3FC894",X"3BCE97",X"2FD397",X"26CB93",X"20B887",X"25C98A",X"2DBD88",X"2EB187",X"40C79C",X"2FC691",X"2FD397",X"17C98B",X"0BC78A",X"00D48F",X"03C68A",X"0DC98F",X"0BC88E",X"01CD8E",X"09DA98",X"3CC59B",X"354C46",X"120000",X"481856",X"630D7A",X"751778",X"320639",X"01061C",X"1D0421",X"7E234F",X"A90D5E",X"C20F73",X"C3006B",X"C20060",X"CD0871",X"C70679",X"B40973",X"B11F72",X"6B3A40",X"2F0C13",X"160309",X"1C1618",X"000300",X"1D3623",X"205133",X"165A35",X"055719",X"0B5520",X"1A5D32",X"276840",X"12572A",X"0A5423",X"0F5D2B",X"0A5929",X"135E33",X"146C3C",X"0B6130",X"1B6333",X"006429",X"07612E",X"1E7940",X"006721",X"157536",X"0B642A",X"175935",X"001D1B",X"0F001D",X"410A43",X"791E7D",X"8A1597",X"8A0C9C",X"7E0288",X"851486",X"4B004E",X"130015",X"28170D",X"733B16",X"DA6E40",X"ED650D",X"EC5A05",X"F76414",X"ED6211",X"F4690E",X"F76707",X"F06C19",X"D86725",X"441500",X"170600",X"1A1A24",X"706664",X"9F836D",X"A58A6D",X"534930",X"141702",X"0B0000",X"E3DCCA"),
(X"FFFEFF",X"7CC9B9",X"04B48E",X"2ABCA5",X"259484",X"000F14",X"0F000D",X"2C1C29",X"531858",X"5E0E55",X"630857",X"4B004D",X"5D0C68",X"7B117D",X"920C89",X"940488",X"95078D",X"96039A",X"8D0095",X"8C028D",X"96028A",X"9E0091",X"9A0095",X"8D038E",X"7A0F6D",X"370741",X"0E0008",X"5D2800",X"E97F27",X"F97C04",X"F97900",X"FF7C0D",X"F47A0D",X"F37308",X"FE770C",X"FF7504",X"FF7901",X"F87600",X"F88005",X"F28006",X"EE7700",X"F57D05",X"FA7D05",X"FA7800",X"F87201",X"F2740E",X"F07E28",X"F18940",X"D67838",X"C97745",X"B67758",X"744C44",X"120001",X"030005",X"000105",X"091113",X"002221",X"0F3F43",X"164D52",X"0F4C51",X"226669",X"0A5359",X"1B6E74",X"005962",X"005955",X"025C5A",X"025658",X"106164",X"0C5D60",X"07605E",X"00615A",X"006259",X"096162",X"075D5E",X"075B5B",X"0A5F5C",X"0C5E5C",X"085A56",X"0B5D59",X"11635D",X"1A5C5B",X"1D5A5B",X"1F565B",X"204F59",X"1F4753",X"2C4D5C",X"264351",X"24404E",X"254240",X"06090E",X"000300",X"7C0847",X"DA1476",X"E60075",X"E20077",X"E70079",X"E60C96",X"E80885",X"BD0A65",X"F09EC6",X"FDF4F7",X"F6FFFC",X"F9FAFE",X"FAFFFF",X"FDFAFF",X"FFFAF2",X"FFFFEF",X"F2FDF9",X"FFFEFF",X"CCBAB0",X"020204",X"3E6380",X"246BD5",X"0676DA",X"0275D0",X"0C66D4",X"1866E4",X"3060B4",X"112236",X"05110F",X"13000E",X"E3D1DF",X"FFFCFE",X"FFFFFB",X"FFFEFF",X"FAF8FB",X"FFFFFF",X"F9FDFC",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FEFEFE",X"FEFEFE",X"FFFFFF",X"F4F4F4",X"20232C",X"686400",X"E2C543",X"F7D327",X"EDCC1F",X"E5C41F",X"F2CE30",X"E5B81D",X"DDB81F",X"E4C826",X"E4D34F",X"FFFBBA",X"FFFFF4",X"F8FCFB",X"FFFFFD",X"FBF6FA",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FCF7FB",X"FDFDF5",X"FFFEFB",X"FAF4C2",X"D9D540",X"EDE046",X"F7E843",X"E7DA33",X"EAE533",X"EAE027",X"EDDE23",X"ECE51B",X"DCD30A",X"DBD922",X"E3CD18",X"F0ED90",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFFF4",X"FFFEFD",X"FFFDF4",X"FFFCCB",X"D8D43D",X"C9C234",X"A09813",X"615300",X"180100",X"000600",X"0D0A03",X"2C2421",X"070602",X"64264F",X"840D4F",X"C05C7E",X"F5E4EA",X"FFFAFF",X"FBFCFF",X"FCFFFF",X"FDFFFC",X"FFFDFE",X"FFFBFF",X"FEF8FF",X"FFEDFF",X"E16AA4",X"C1035B",X"D81070",X"C80D66",X"A91859",X"44041E",X"000200",X"02603C",X"22956A",X"22A675",X"17A06C",X"23B67F",X"1DC185",X"18BD85",X"13AB7A",X"1ABE7F",X"10A06B",X"189B71",X"27AE83",X"0AA16C",X"14B87C",X"1DCF91",X"10CC8F",X"04DD98",X"07CA8E",X"0ECA90",X"10CD93",X"07D394",X"0BDC9A",X"20A97F",X"000F09",X"150000",X"491957",X"6D1784",X"6D0F70",X"4D2154",X"00041A",X"0F0013",X"6D123E",X"B71B6C",X"D11E82",X"E11D89",X"D20B70",X"CA056E",X"CD0C7F",X"CC218B",X"8B004C",X"2B0000",X"1F0003",X"0D0000",X"040000",X"121912",X"0E2714",X"1F5032",X"20643F",X"0E6022",X"155F2A",X"1F6237",X"25663E",X"02471A",X"1C6635",X"277543",X"156434",X"236E43",X"015929",X"095F2E",X"236B3B",X"016A2F",X"045E2B",X"0A652C",X"006620",X"046425",X"0C652B",X"003D19",X"000F0D",X"070015",X"420B44",X"680D6C",X"760183",X"840696",X"73007D",X"811082",X"5B0E5E",X"280B2A",X"190800",X"68300B",X"B64A1C",X"F36B13",X"F6640F",X"F66313",X"EF6413",X"EA5F04",X"FF6F0F",X"E25E0B",X"E77634",X"895A3C",X"0D0000",X"000009",X"6F6563",X"997D67",X"63482B",X"2B2108",X"010400",X"201400",X"DED7C5"),
(X"FEFFFD",X"8BABA6",X"1AA584",X"2FAE93",X"16584E",X"000408",X"000807",X"00150D",X"001900",X"001100",X"000F00",X"001200",X"00120B",X"000515",X"300C30",X"430C36",X"691D77",X"891091",X"920094",X"920092",X"920794",X"900197",X"900499",X"870790",X"83037A",X"3C074F",X"07000A",X"521D00",X"E97A33",X"FF841E",X"FF7E09",X"FA7703",X"FF730F",X"FF6B07",X"FF710A",X"FF7506",X"FF7B05",X"FC7800",X"FF7C05",X"FF7A07",X"F77500",X"F97705",X"F97509",X"FD740A",X"FF7B0C",X"FF7902",X"F87400",X"F07300",X"FF7B19",X"FF801B",X"F77D18",X"E07316",X"B95D10",X"974B17",X"440700",X"270000",X"150000",X"0D0000",X"0A0905",X"202F2C",X"122C29",X"153C39",X"2D5D5F",X"356C71",X"0B555E",X"0D5C63",X"02555B",X"065E62",X"005556",X"005655",X"065854",X"0C5B56",X"155B5D",X"0C5A5A",X"055E5A",X"04655E",X"04655E",X"055E5A",X"0B5A57",X"145A5A",X"00605F",X"005D5C",X"005B5D",X"045D61",X"045E5F",X"0D6768",X"076161",X"0A6663",X"295E58",X"112027",X"000A00",X"700D4D",X"CA1974",X"DF0575",X"DA057B",X"D5007E",X"C40576",X"CA2A84",X"86134E",X"CC87A6",X"FFF4FF",X"FDFBFE",X"F7FBFC",X"FFFFFF",X"F5FCF4",X"FFFCFD",X"FFF6FF",X"F9FFFF",X"FAFEFF",X"E7E4ED",X"4961A1",X"165CD6",X"0B6EE3",X"0B6AE0",X"0669E8",X"107DF2",X"0075DF",X"006EE7",X"1151BD",X"21265D",X"000014",X"A29EAD",X"FFFCFF",X"FAF6F7",X"F6F8F7",X"F7FBFC",X"FEFFFF",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FEFEFE",X"FEFEFE",X"FFFFFF",X"F4F4F4",X"292D30",X"424122",X"9A8A71",X"A58E62",X"99815F",X"938055",X"AB9B79",X"AD9F78",X"AC8870",X"AD8E71",X"9F8971",X"F9EFE6",X"FDFDFF",X"F6FAFD",X"FFFFFD",X"FFFDFA",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"F7FEEE",X"FEFEF6",X"FDF3AE",X"E5D810",X"F0D313",X"ECD00A",X"F4DF14",X"ECDD06",X"EEDE05",X"E7CF00",X"F0E309",X"EEDF08",X"DFDB18",X"F8D40C",X"F5F2A1",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"F2F9FF",X"FBFFFF",X"F3F7F6",X"F8F8FF",X"C9CDB2",X"010500",X"040100",X"050000",X"0A0200",X"2C3500",X"74742E",X"3E3E1A",X"040000",X"6F2854",X"B52F76",X"92132E",X"EED1ED",X"FFF9FF",X"F5F4F9",X"FAFEFD",X"FFFFFF",X"FFFCFD",X"FAF8FB",X"FBFCFE",X"F6FDFF",X"F7B7D9",X"A1074F",X"DD1673",X"C70464",X"B61160",X"5F0028",X"1B0006",X"0E0002",X"08050C",X"00040A",X"0E151B",X"162425",X"274640",X"203F3A",X"3F5354",X"12050E",X"201A24",X"16232B",X"1A2E2F",X"000908",X"000A00",X"29926A",X"0ED18D",X"0DCD91",X"11C48C",X"13C68E",X"0DCA90",X"00CB8C",X"0BD697",X"209E79",X"000305",X"0C1019",X"40184C",X"7D2780",X"80217D",X"6D216C",X"3E0844",X"1D0022",X"2E0D2A",X"5C1734",X"B1297B",X"D4148D",X"C20070",X"B11463",X"972C60",X"481D2E",X"12180A",X"1F040B",X"1A1200",X"AEB936",X"8F9720",X"0B0500",X"1B1217",X"101C1A",X"1D3F1E",X"225149",X"2E6457",X"2C705B",X"09633D",X"00632A",X"006F2F",X"0D7334",X"0B642C",X"137334",X"005E1B",X"006322",X"1C6B3C",X"096F3F",X"0F5D35",X"0B5D2F",X"0C5E30",X"20503A",X"386048",X"051717",X"10012C",X"37014C",X"630661",X"820C7C",X"7D0083",X"7C0096",X"8523AA",X"6F1189",X"760878",X"5A0057",X"1F0025",X"2A0D21",X"3A0B13",X"BF582D",X"F07C33",X"E16004",X"F3660E",X"F95A08",X"FF5C06",X"F9680B",X"EE781E",X"CC6731",X"400700",X"0D0009",X"463B4B",X"5B504E",X"171000",X"0A0200",X"52460C",X"9D912D",X"F9F298"),
(X"FCFEFB",X"7C9C97",X"079271",X"2FAE93",X"00342A",X"000307",X"192D2C",X"2B544C",X"32785E",X"497A65",X"4A7561",X"447967",X"39645D",X"101626",X"150015",X"2C001F",X"540862",X"850C8D",X"940096",X"930093",X"8F0491",X"8C0093",X"91059A",X"8B0B94",X"8A0A81",X"3B064E",X"060009",X"562101",X"E1722B",X"FF851F",X"FF800B",X"F97602",X"FF7511",X"FF6B07",X"FF710A",X"FF7708",X"FF7E08",X"FD7900",X"FF7D06",X"FF7C09",X"FE7C04",X"F97705",X"F36F03",X"F56C02",X"FB6F00",X"FB7000",X"FA7600",X"FD8000",X"F46A08",X"F36F0A",X"F47A15",X"F38629",X"E28639",X"D88C58",X"A5684B",X"885345",X"866A5F",X"180700",X"010000",X"000A07",X"000D0A",X"001B18",X"063638",X"00363B",X"0E5861",X"0F5E65",X"085B61",X"086064",X"025A5B",X"015756",X"095B57",X"0E5D58",X"145A5C",X"0A5858",X"005955",X"005D56",X"005F58",X"035C58",X"0B5A57",X"125858",X"026463",X"016160",X"036163",X"0A6367",X"035D5E",X"066061",X"045E5E",X"0F6B68",X"285D57",X"1F2E35",X"000C00",X"630040",X"C5146F",X"DE0474",X"D60177",X"DA0583",X"D21384",X"9C0056",X"590021",X"601B3A",X"F7DBE9",X"FEFCFF",X"F8FCFD",X"FBFBFD",X"FBFFFA",X"FFFCFD",X"FFF4FF",X"F3F9FF",X"F3F7FA",X"F9F6FF",X"859DDD",X"0E54CE",X"1376EB",X"0968DE",X"076AE9",X"0976EB",X"0176E0",X"0270E9",X"2D6DD9",X"292E65",X"000014",X"221E2D",X"EEE7EE",X"FFFEFF",X"FEFFFF",X"FBFFFF",X"FDFEFF",X"FEFCFD",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FEFEFE",X"FEFEFE",X"FFFFFF",X"F4F4F4",X"393D40",X"040300",X"140400",X"150000",X"150000",X"130000",X"110100",X"0E0000",X"1F0000",X"1C0000",X"120000",X"EAE0D7",X"FFFFFF",X"FCFFFF",X"F8F8F6",X"FFFEFB",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FCFDFF",X"F8FFEF",X"FFFFF8",X"FBF1AC",X"E2D50D",X"F5D818",X"E8CC06",X"F5E015",X"E9DA03",X"EADA01",X"F1D907",X"E5D800",X"E8D902",X"E4E01D",X"EFCB03",X"FBF8A7",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"F8FFFF",X"F9FFFD",X"FCFFFF",X"F9F9FF",X"CDD1B6",X"040800",X"2B2823",X"342F2B",X"938B64",X"C4CD7A",X"DBDB95",X"6F6F4B",X"040000",X"510A36",X"A21C63",X"71000D",X"A98CA8",X"FFF7FF",X"FFFEFF",X"F3F7F6",X"FAFAFA",X"FFFEFF",X"FFFEFF",X"F7F8FA",X"F8FFFF",X"FFD4F6",X"C52B73",X"CB0461",X"D41171",X"B40F5E",X"7A1243",X"320B1D",X"1B060F",X"08050C",X"000208",X"000107",X"000506",X"001711",X"000A05",X"000F10",X"0C0008",X"0D0711",X"00060E",X"000A0B",X"0A1312",X"000900",X"137C54",X"07CA86",X"00C084",X"0DC088",X"11C48C",X"0ECB91",X"00CA8B",X"08D394",X"1C9A75",X"000305",X"11151E",X"23002F",X"5C065F",X"8B2C88",X"5C105B",X"5B2561",X"27002C",X"170013",X"37000F",X"90085A",X"CC0C85",X"CD0B7B",X"BA1D6C",X"6D0236",X"2D0213",X"000500",X"3C2128",X"ADA564",X"C5D04D",X"CED65F",X"7A7442",X"0B0207",X"000B09",X"072908",X"0D3C34",X"174D40",X"226651",X"1A744E",X"00682F",X"006D2D",X"006627",X"09622A",X"127233",X"137431",X"005B1A",X"105F30",X"0E7444",X"1C6A42",X"1F7143",X"06582A",X"093923",X"052D15",X"000A0A",X"060022",X"450F5A",X"741772",X"7F0979",X"87038D",X"7E0098",X"741299",X"761890",X"7C0E7E",X"741571",X"3E0D44",X"1D0014",X"200000",X"AD461B",X"EB772E",X"ED6C10",X"EA5D05",X"FE5F0D",X"FF5B05",X"F9680B",X"DF690F",X"DB7640",X"713827",X"12000E",X"2A1F2F",X"0E0301",X"181100",X"4C441D",X"9D9157",X"AB9F3B",X"E6DF85"),
(X"F4FEF6",X"A88A96",X"195748",X"4F8D80",X"060A0D",X"000A04",X"16936B",X"2DE0A8",X"1BD4B2",X"2BDFB8",X"1BD9A9",X"18E5AD",X"32E8B8",X"26997C",X"00251B",X"000000",X"2B052E",X"790D70",X"9F008F",X"9A0094",X"8B0598",X"850098",X"98019E",X"A00094",X"701783",X"220B39",X"060500",X"7D4401",X"EC7316",X"FF7E0B",X"F97C00",X"FB7F00",X"FC8100",X"EF7800",X"F18000",X"F38700",X"F68A04",X"F17F05",X"FB8018",X"FE7F22",X"F97513",X"F07112",X"EE7313",X"F57B16",X"F87910",X"F66F03",X"FA6F06",X"FF7912",X"FC860B",X"F57900",X"FC7A00",X"FB7802",X"E36D03",X"E28029",X"DA9049",X"C68950",X"C19169",X"865938",X"5D381E",X"563320",X"170000",X"110000",X"0A0000",X"060201",X"1E201D",X"222C2B",X"233D3C",X"275052",X"265D60",X"165A5D",X"10595F",X"075257",X"006059",X"005F5B",X"055D5E",X"095C60",X"0C5F65",X"096067",X"016066",X"005C60",X"025A5C",X"03585B",X"08595D",X"0B5A5F",X"035256",X"075758",X"055755",X"126460",X"14535C",X"151433",X"080000",X"6F0550",X"CB1D76",X"E7046F",X"E40074",X"E30282",X"D20D5F",X"580027",X"18171D",X"000708",X"BCBFC4",X"F4FEFF",X"F7FDFB",X"FFFBF9",X"F0FEFE",X"FFF9FF",X"FFF9FF",X"F8FDF9",X"FCFFF1",X"FBFFFC",X"99C6F0",X"046CC5",X"1D7BD3",X"0074E1",X"097EF0",X"096BD6",X"006CD6",X"0173E5",X"0F6FDF",X"005AC1",X"102A3B",X"000410",X"C9C8CE",X"FFFEFF",X"F2F8F6",X"F3FCFB",X"FFFFFF",X"FFFBFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FEFEFE",X"FEFEFE",X"FFFFFF",X"F4F4F4",X"3A3728",X"080000",X"2E1421",X"2A0200",X"38000A",X"3C0000",X"350000",X"3B0100",X"190200",X"28140D",X"0B0000",X"ECE8DD",X"F7FAF3",X"FCFFFF",X"FDFCFF",X"FFFDFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FBFCFF",X"F7FFF8",X"FDFEF8",X"F2EAA1",X"E0D500",X"FCE118",X"EEDA07",X"E6DD02",X"EED904",X"F1DC09",X"ECCF09",X"E6D607",X"F2DE0E",X"E8E01D",X"FCCF00",X"EEE995",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFAFD",X"FFFDF2",X"FEFBF2",X"FFFFFD",X"EAE6F7",X"6B6766",X"04000C",X"9B9C63",X"EDF473",X"E7E926",X"DDDB2E",X"757B31",X"000600",X"1E1216",X"1B0005",X"230209",X"2A0B11",X"E1D2CF",X"FFFFF6",X"FDFFFA",X"F7F6FC",X"FFFBFF",X"FEFEFF",X"F9FEF7",X"FBFFFC",X"FCF3F8",X"DB8AB3",X"AA085B",X"D7147D",X"CB006E",X"C20D6E",X"8F0D55",X"9C0046",X"8F034C",X"930F5B",X"950655",X"A10D59",X"9E1058",X"9A0E55",X"91004A",X"8E1059",X"9E065B",X"AB166A",X"851658",X"632049",X"150414",X"145D4A",X"24C695",X"0BCF8F",X"01CC8A",X"00CD88",X"02DB97",X"07D998",X"0AD89A",X"06996F",X"001107",X"0A1318",X"000402",X"0A1511",X"110F1A",X"1B0124",X"44184D",X"451D51",X"130022",X"050215",X"510F3F",X"8F285F",X"732D47",X"1E0B05",X"343219",X"0D0400",X"605000",X"C4B011",X"E5DB2E",X"CFCE11",X"E9E222",X"D7C71A",X"C2AF2F",X"453D00",X"020700",X"222826",X"152822",X"193E2D",X"346649",X"124A25",X"225C36",X"1A5535",X"236247",X"115C31",X"256B39",X"0C602C",X"1F5A3A",X"145B39",X"1D4125",X"224531",X"1A292E",X"0E011F",X"0A0012",X"280837",X"3F0A62",X"5E0E81",X"7E128A",X"7D0483",X"9015A3",X"8B1A84",X"A72B9D",X"7B037E",X"6D0985",X"8F30A8",X"660B6B",X"260026",X"000606",X"663E34",X"CA6B33",X"FF7518",X"F25100",X"F25909",X"FB6913",X"F76404",X"F66701",X"FD6E12",X"B95D2A",X"250000",X"090000",X"000300",X"353F1C",X"9D9648",X"D0AD39",X"B69F2D",X"F7E47E"),
(X"F9FFFB",X"A58793",X"001405",X"155346",X"000104",X"172A24",X"3EBB93",X"1ED199",X"15CEAC",X"1ACEA7",X"16D4A4",X"09D69E",X"24DAAA",X"53C6A9",X"285248",X"000000",X"250028",X"780C6F",X"A00090",X"9D0097",X"900A9D",X"8B049E",X"9B04A1",X"9E0092",X"69107C",X"16002D",X"0B0A00",X"9D6421",X"FA8124",X"FF800D",X"F77A00",X"FF8300",X"FC8100",X"F07900",X"F48300",X"F68A03",X"F88C06",X"F17F05",X"FB8018",X"FF8225",X"FF811F",X"FF8223",X"FE8323",X"F87E19",X"F17209",X"F66F03",X"FF740B",X"FF7710",X"F98308",X"FB7F03",X"F87600",X"FC7903",X"F98319",X"D5731C",X"9C520B",X"6D3000",X"693911",X"663918",X"59341A",X"A5826F",X"8C6F61",X"301A0F",X"090000",X"040000",X"020401",X"000807",X"001615",X"022B2D",X"11484B",X"0D5154",X"155E64",X"0F5A5F",X"00645D",X"03635F",X"055D5E",X"04575B",X"05585E",X"075E65",X"026167",X"005F63",X"065E60",X"075C5F",X"095A5E",X"0B5A5F",X"065559",X"0D5D5E",X"095B59",X"11635F",X"195861",X"0A0928",X"090000",X"7D135E",X"C61871",X"E3006B",X"EB037B",X"DD007C",X"D40F61",X"721541",X"0B0A10",X"000405",X"888B90",X"F2FCFE",X"FBFFFF",X"FFF6F4",X"F2FFFF",X"FFFBFF",X"FFF3FD",X"FAFFFB",X"FCFFF1",X"F7FCF8",X"D0FDFF",X"0B73CC",X"1371C9",X"017BE8",X"0277E9",X"0E70DB",X"006FD9",X"0375E7",X"0969D9",X"1672D9",X"3B5566",X"00020E",X"7C7B81",X"FEFCFD",X"FAFFFE",X"F9FFFF",X"FCFCFC",X"FFFAFE",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FEFEFE",X"FEFEFE",X"FFFFFF",X"F4F4F4",X"3D3A2B",X"0A0000",X"3A202D",X"3D1513",X"541A26",X"5A1B12",X"46080B",X"4B110F",X"3A231B",X"37231C",X"0B0000",X"E8E4D9",X"FEFFFA",X"FBFFFF",X"FFFEFF",X"FEF9FF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FCFDFF",X"F7FFF8",X"FFFFFA",X"FFF7AE",X"E7DC04",X"EFD40B",X"ECD805",X"E9E005",X"EFDA05",X"E9D401",X"F2D50F",X"E6D607",X"EAD606",X"E4DC19",X"FCCF00",X"FBF6A2",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFAFD",X"FFFFF4",X"FFFCF3",X"FFFEFC",X"FFFCFF",X"938F8E",X"090011",X"616229",X"CFD655",X"E8EA27",X"DAD82B",X"61671D",X"000500",X"1F1317",X"3D1C27",X"35141B",X"150000",X"CBBCB9",X"F8F8EE",X"FAFCF7",X"FFFEFF",X"FFFCFF",X"FBFBFD",X"FCFFFA",X"FAFFFB",X"FFFCFF",X"FFBCE5",X"BC1A6D",X"C4016A",X"D10574",X"BE096A",X"A5236B",X"BB1B65",X"AD216A",X"9B1763",X"B62776",X"AC1864",X"AC1E66",X"AF236A",X"B01E69",X"A2246D",X"AF176C",X"B52074",X"A63779",X"6F2C55",X"0A0009",X"19624F",X"1DBF8E",X"0BCF8F",X"04CF8D",X"00CE89",X"00D793",X"00D08F",X"0DDB9D",X"36C99F",X"3C7167",X"020B10",X"000503",X"000400",X"01000A",X"0F0018",X"25002E",X"3B1347",X"341B43",X"020012",X"4C0A3A",X"750E45",X"440018",X"0E0000",X"0D0B00",X"B0A76E",X"DBCB73",X"EDD93A",X"D2C81B",X"D4D316",X"D1CA0A",X"E9D92C",X"E8D555",X"C2BA6F",X"565B32",X"060C0A",X"000600",X"000D00",X"002306",X"003813",X"104A24",X"114C2C",X"2C6B50",X"206B40",X"185E2C",X"085C28",X"104B2B",X"003917",X"001700",X"001200",X"041318",X"120523",X"1B0923",X"2C0C3B",X"7A459D",X"7B2B9E",X"7D1189",X"8C1392",X"7D0290",X"84137D",X"A32799",X"750078",X"85219D",X"771890",X"7A1F7F",X"401240",X"000808",X"1D0000",X"AF5018",X"FF6C0F",X"FF6308",X"F25909",X"F4620C",X"F76404",X"F46500",X"FD6E12",X"BA5E2B",X"2C0600",X"221819",X"000300",X"6F7956",X"B1AA5C",X"C7A430",X"C1AA38",X"FFEF89"),
(X"F8FFFF",X"AB8B9A",X"000800",X"272121",X"010204",X"0A7D5C",X"2DE4AC",X"03DA96",X"00D59F",X"09DDA0",X"0BE79F",X"03D999",X"16E2AD",X"20E2B0",X"006A48",X"070000",X"2B0A27",X"700C6C",X"980792",X"8C008C",X"92048A",X"A00295",X"93058B",X"7C1683",X"3D1039",X"160002",X"390700",X"C56721",X"FF881A",X"FF8704",X"FC7500",X"FF7C0F",X"F5810A",X"FB8300",X"FF8100",X"F67309",X"F78129",X"E17946",X"CE6A5B",X"B14C40",X"9D6F62",X"946E5B",X"845F33",X"95612F",X"D88B43",X"F18336",X"F47025",X"F37800",X"FF7803",X"EA750C",X"F47A24",X"F5853D",X"B17C48",X"332518",X"04000C",X"000013",X"000A28",X"000017",X"000110",X"40292F",X"977C6B",X"BB8757",X"C66521",X"844500",X"1C0000",X"180000",X"190000",X"120000",X"0A0000",X"080A07",X"172727",X"23383B",X"264C59",X"245462",X"1D5866",X"145A62",X"105A5D",X"0B5753",X"065751",X"095B57",X"0D6356",X"066054",X"015E54",X"005E57",X"005B57",X"005A59",X"045C5D",X"0C5F63",X"124F52",X"181F27",X"0E0001",X"75103C",X"D81476",X"D70077",X"DF0080",X"E0047F",X"D30975",X"B30F66",X"5A0033",X"0B000A",X"63746E",X"E6ECEA",X"FDFCFF",X"F5FAFF",X"FFFAFF",X"FFFDFF",X"FFFFFD",X"FFFFFA",X"FDFCFA",X"FCFFFF",X"EFFBFF",X"98ABBA",X"0660D8",X"1D72E7",X"1976EF",X"0066E6",X"0776EC",X"0469D3",X"046BD0",X"0373E1",X"1667DA",X"002569",X"000010",X"DBD1D0",X"FFFEFF",X"FBF6FC",X"FFFAFD",X"FFFDFB",X"FCFFFF",X"FFFFFF",X"FFFEFC",X"FFFFFD",X"FCFFFF",X"FBFFFF",X"FEFEFF",X"F6F2F1",X"2F3533",X"090305",X"7E1E39",X"C00F3D",X"BC0E31",X"C31435",X"C1092F",X"B61235",X"A42341",X"57141B",X"0B0200",X"E0E9D6",X"FFFFFD",X"FFF6FF",X"FFFCFF",X"F6FEF1",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFDFF",X"FCF8F5",X"F2FFEA",X"F2F1B8",X"DACD71",X"EED861",X"FAE160",X"E2EB5C",X"EEE25A",X"EFDD33",X"F6E758",X"FBD832",X"EBD544",X"E7EC5E",X"E4DA2A",X"FAF0BF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FEFEFE",X"FFFFFD",X"F9F7FF",X"FFFFF8",X"DFDBDA",X"040000",X"6E7A00",X"DCE944",X"EAE71C",X"E5DA33",X"7A7821",X"0A0000",X"491C19",X"6E1727",X"861B39",X"5A0006",X"B65868",X"FFE5E9",X"FFFBF9",X"FEFEFC",X"FFFCFF",X"FFF6FF",X"F7FFFF",X"FFFAF8",X"FBFFFB",X"FFEEF6",X"CD759F",X"A60352",X"D61777",X"C50E6B",X"B30962",X"BF0A71",X"CC0071",X"DC097E",X"B2066C",X"C61275",X"D0036A",X"C6086A",X"CD006B",X"CB0478",X"CD0474",X"D60068",X"DC207E",X"80285B",X"02020E",X"1A5745",X"4ABF93",X"1AC893",X"1BCC95",X"1FC690",X"19B681",X"19C88F",X"19DB9E",X"1EC693",X"3DB494",X"229878",X"2D9E80",X"06735C",X"104E4B",X"003428",X"000306",X"381943",X"5A116D",X"24004B",X"260939",X"1C0110",X"110000",X"353511",X"9A9E4A",X"D2D13B",X"DEDD13",X"E5D000",X"E8D00E",X"E7CA16",X"E4C709",X"E7CE02",X"DAC810",X"E3D453",X"DDD282",X"33392B",X"000300",X"0F1312",X"050304",X"120000",X"1A0804",X"162413",X"0D180A",X"2B3E3C",X"14292A",X"00000C",X"110010",X"1D0012",X"1F001D",X"180022",X"320240",X"480264",X"611378",X"59006A",X"9535A3",X"A23EB0",X"821B8E",X"84178E",X"75037C",X"660681",X"790284",X"790078",X"962496",X"8C1D96",X"8A1A98",X"7A247D",X"2D0025",X"070001",X"7E462D",X"EE7A3D",X"FD6512",X"F45900",X"F9650D",X"F06007",X"FA690C",X"F05802",X"D7712F",X"7F492D",X"0A0001",X"0E0112",X"294A43",X"505F4A",X"8E6F5A",X"9D915D",X"FCEEC9"),
(X"F8FFFF",X"AE8E9D",X"000B02",X"2C2626",X"000002",X"2DA07F",X"26DDA5",X"0AE19D",X"08DEA8",X"06DA9D",X"08E49C",X"02D898",X"0EDAA5",X"23E5B3",X"1A8C6A",X"0A0100",X"2E0D2A",X"771373",X"94038E",X"920592",X"96088E",X"9C0091",X"95078D",X"710B78",X"290025",X"180004",X"744229",X"E3853F",X"FF8113",X"FF7B00",X"FF7B00",X"FF780B",X"F37F08",X"FA8200",X"FF8201",X"FE7B11",X"ED771F",X"AC4411",X"570000",X"660100",X"220000",X"1D0000",X"240000",X"2A0000",X"8D4000",X"D6681B",X"F67227",X"FF8604",X"FF7300",X"F07B12",X"F47A24",X"D6661E",X"350000",X"0B0000",X"0F0617",X"1B2034",X"1A3553",X"2C344B",X"141625",X"100000",X"1B0000",X"9A6636",X"FC9B57",X"C58636",X"8D7050",X"725438",X"573D26",X"2E180A",X"0B0100",X"000100",X"000808",X"000B0E",X"00202D",X"073745",X"0F4A58",X"0F555D",X"166063",X"1A6662",X"12635D",X"0B5D59",X"065C4F",X"035D51",X"036056",X"02635C",X"01615D",X"015D5C",X"025A5B",X"075A5E",X"165356",X"10171F",X"0E0001",X"77123E",X"D91577",X"DE027E",X"E10082",X"DF037E",X"D80E7A",X"BE1A71",X"71174A",X"0D000C",X"000C06",X"B6BCBA",X"F9F8FD",X"FBFFFF",X"FFFBFF",X"FDFBFE",X"FEFEFC",X"FFFEF9",X"FFFFFD",X"FBFEFF",X"F4FFFF",X"C6D9E8",X"0660D8",X"166BE0",X"0E6BE4",X"127DFD",X"006DE3",X"0D72DC",X"056CD1",X"0373E1",X"1465D8",X"294E92",X"090619",X"A79D9C",X"FFFEFF",X"FFFDFF",X"FFFCFF",X"FFFAF8",X"FCFFFF",X"FFFFFF",X"FFFEFC",X"FFFFFD",X"FCFFFF",X"FBFFFF",X"FEFEFF",X"F6F2F1",X"363C3A",X"040000",X"7B1B36",X"B80735",X"BD0F32",X"B70829",X"BF072D",X"B51134",X"971634",X"49060D",X"080000",X"E2EBD8",X"FFFFFD",X"FFF5FF",X"FFFCFF",X"FBFFF6",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FCF7FB",X"FFFEFB",X"F2FFEA",X"C9C88F",X"554800",X"846E00",X"A78E0D",X"9BA415",X"B5A921",X"BBA900",X"BCAD1E",X"E5C21C",X"C6B01F",X"B7BC2E",X"A39900",X"DAD09F",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FBFBFB",X"FFFFFD",X"FEFCFF",X"FFFFF7",X"F9F5F4",X"5F5B52",X"889416",X"E0ED48",X"E8E51A",X"F8ED46",X"A2A049",X"080000",X"512421",X"761F2F",X"740927",X"83232F",X"6D0F1F",X"E8BEC2",X"FFF6F4",X"FDFDFB",X"FFFBFF",X"FFF8FF",X"F0FBFF",X"FFF9F7",X"F8FFF8",X"FFF6FE",X"FFB2DC",X"A80554",X"D01171",X"C20B68",X"C0166F",X"BE0970",X"D10576",X"DE0B80",X"BC1076",X"C91578",X"CF0269",X"C50769",X"D1036F",X"C50072",X"C90070",X"D70069",X"CE1270",X"660E41",X"00000B",X"1D5A48",X"44B98D",X"18C691",X"0DBE87",X"24CB95",X"2DCA95",X"1BCA91",X"1ADC9F",X"25CD9A",X"30A787",X"41B797",X"47B89A",X"50BDA6",X"6EACA9",X"2C6E62",X"000407",X"2C0D37",X"681F7B",X"441E6B",X"110024",X"230817",X"0E0000",X"3E3E1A",X"CBCF7B",X"DEDD47",X"CFCE04",X"E8D300",X"E4CC0A",X"E9CC18",X"EDD012",X"DBC200",X"F5E32B",X"D5C645",X"8C8131",X"000300",X"0F120B",X"030706",X"232122",X"280D12",X"140200",X"000600",X"000500",X"000604",X"000F10",X"00020E",X"381B37",X"441539",X"390C37",X"461B50",X"3C0C4A",X"561072",X"6A1C81",X"670E78",X"71117F",X"6C087A",X"61006D",X"8B1E95",X"86148D",X"8626A1",X"AC35B7",X"7E007D",X"710071",X"6F0079",X"740482",X"77217A",X"47173F",X"060000",X"7C442B",X"DF6B2E",X"FE6613",X"FD6208",X"FF6D15",X"FE6E15",X"EA5900",X"FF6812",X"DD7735",X"804A2E",X"0F0506",X"241728",X"12332C",X"000C00",X"180000",X"120600",X"D6C8A3"),
(X"FFFAFF",X"B38D9C",X"000500",X"121210",X"004428",X"36D2A3",X"00E19B",X"08DF9B",X"08EEA5",X"00DC8F",X"00E792",X"00E893",X"13DE9C",X"3FD2A8",X"216556",X"060004",X"41054F",X"84158B",X"92009F",X"9A089B",X"9A059F",X"960087",X"851384",X"491152",X"060011",X"421300",X"CD6E1C",X"FF8B10",X"FA8501",X"EF7F02",X"F1820C",X"F07F09",X"FF7C15",X"FF8A05",X"F67E10",X"DC874E",X"865E3B",X"0F0000",X"180420",X"180035",X"35002E",X"350031",X"260020",X"27002C",X"140007",X"240900",X"A77763",X"D08238",X"E37F05",X"FF9013",X"D47839",X"370A0F",X"0E0014",X"101646",X"1C47A6",X"1C66D3",X"1471DB",X"1966DA",X"215DBD",X"001750",X"000007",X"340A00",X"CF7340",X"EB9528",X"FE8A13",X"F48212",X"F28624",X"D77828",X"904106",X"4B0F00",X"220000",X"190000",X"000400",X"050C00",X"07100B",X"0A1415",X"142223",X"213536",X"264645",X"295150",X"285666",X"265766",X"215966",X"1D5964",X"15555E",X"105359",X"115759",X"155B5B",X"1A4F57",X"05121B",X"060007",X"761149",X"E01183",X"EF0088",X"EE007D",X"E40270",X"DE0882",X"D70978",X"AE1768",X"3C0628",X"000305",X"677872",X"F0F6F2",X"FBFFFA",X"FFFDFF",X"FDFDFF",X"FFFFFD",X"FDFCF8",X"FFFEFF",X"FCFBFF",X"F7FFFF",X"EDFBFF",X"6395C8",X"1362BE",X"117BF3",X"0F7CF1",X"0D77DD",X"0772DA",X"0972E8",X"0667EA",X"066AD9",X"186DDA",X"002C82",X"2F3662",X"EDE4F5",X"F9FBFF",X"F4FDFF",X"FBFFFF",X"FDFEFF",X"FFFFFF",X"FFFEFA",X"FFFFFD",X"FBFFFF",X"FBFFFF",X"FDFEFF",X"F4F3F1",X"403B38",X"070000",X"7E0E24",X"CE012C",X"CF0324",X"C9001C",X"C80023",X"B2132F",X"5B1329",X"15010A",X"0A0102",X"EDE0D8",X"FEFFFA",X"F8F8FF",X"FEF4FD",X"FCFFF6",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFCFF",X"FBEEFF",X"F8FEFF",X"D0CFD5",X"120000",X"130000",X"1C0000",X"1E000D",X"0B0000",X"0D0000",X"120005",X"250001",X"000500",X"2B1A22",X"000300",X"C8BEBC",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"F9F9F9",X"FCFCFA",X"FFFEFF",X"F6F6EE",X"FFFEFF",X"C0BBB8",X"99A239",X"DEE535",X"D3CC02",X"FDF344",X"979E2A",X"130D00",X"4A142B",X"7D0936",X"9D072A",X"921D25",X"67000C",X"CF718B",X"FFEFFB",X"F9FFFF",X"FAFCFB",X"F7FFFF",X"FBFFFF",X"FBFFFF",X"FFFEFF",X"FCF6F8",X"FFF7FF",X"9C6E8A",X"61103B",X"872E5A",X"671B3F",X"6D2040",X"7F244F",X"8D1B56",X"871F5A",X"8A1E5C",X"7D1353",X"80175C",X"B0116D",X"BD1060",X"C50A63",X"CD0568",X"C51373",X"6C0348",X"140013",X"1C302E",X"255D40",X"2F5345",X"143D2D",X"3B6456",X"54756A",X"335C4E",X"336959",X"366C5C",X"0F3D30",X"1C4E43",X"2D5D51",X"2FB995",X"2DBD9A",X"176450",X"090307",X"37153A",X"78086A",X"6F1078",X"490050",X"35003E",X"20042C",X"030000",X"8E8D54",X"DFD454",X"D5C00F",X"E7D51D",X"DBD408",X"D0D500",X"C9D004",X"DDDA3F",X"C1B75E",X"766D4E",X"030000",X"001118",X"1A1826",X"080705",X"5F3A1D",X"B65F29",X"963E00",X"7E3814",X"541714",X"00060B",X"190329",X"470A5A",X"5D0F7C",X"6B118C",X"760E8B",X"6A057D",X"812798",X"942DA0",X"75087D",X"740078",X"850D89",X"8E1893",X"74007B",X"8C1593",X"840986",X"781582",X"AA3FB3",X"872191",X"872594",X"9124A1",X"861195",X"721878",X"320232",X"0C1011",X"906449",X"D1692A",X"F0630B",X"EF5B00",X"F66A08",X"F46A07",X"F86A04",X"EF5D07",X"E46619",X"843B08",X"000100",X"29266B",X"2F41A3",X"13297F",X"12306C",X"00002B",X"D2D7F4"),
(X"FFFAFF",X"B791A0",X"000500",X"000000",X"2B8B6F",X"3BD7A8",X"00DC96",X"09E09C",X"00E59C",X"04E295",X"00E994",X"00E691",X"1CE7A5",X"37CAA0",X"002A1B",X"090007",X"490D57",X"86178D",X"9400A1",X"99079A",X"98039D",X"99018A",X"7B097A",X"390142",X"03000E",X"6B3C22",X"DD7E2C",X"F37D02",X"FF8B07",X"F48407",X"EB7C06",X"F07F09",X"FB760F",X"F97300",X"FF8B1D",X"BF6A31",X"260000",X"0F0000",X"13001B",X"250842",X"501B49",X"551851",X"51184B",X"320637",X"200113",X"1E0300",X"2D0000",X"C4762C",X"F18D13",X"F88609",X"AA4E0F",X"1F0000",X"0E0014",X"343A6A",X"436ECD",X"2872DF",X"116ED8",X"2471E5",X"2E6ACA",X"2A4982",X"0D0D15",X"200000",X"9A3E0B",X"E79124",X"F6820B",X"F38111",X"F18523",X"EA8B3B",X"D5864B",X"C28661",X"865942",X"4E2D1E",X"010500",X"000600",X"000702",X"040E0F",X"031112",X"000B0C",X"000A09",X"000F0E",X"0A3848",X"0F404F",X"144C59",X"17535E",X"16565F",X"16595F",X"1C6264",X"226868",X"164B53",X"0E1B24",X"060007",X"710C44",X"DE0F81",X"E90082",X"EE007D",X"E70573",X"D8027C",X"D40675",X"B72071",X"541E40",X"091416",X"000E08",X"C1C7C3",X"F9FEF8",X"FCFAFF",X"FCFCFE",X"FFFFFD",X"FFFEFA",X"FFFDFE",X"FFFEFF",X"F6FFFF",X"F2FFFF",X"94C6F9",X"0958B4",X"0872EA",X"0976EB",X"0973D9",X"0974DC",X"046DE3",X"0C6DF0",X"0C70DF",X"176CD9",X"2B59AF",X"000430",X"B8AFC0",X"FCFEFF",X"F1FAFF",X"FBFFFF",X"FDFEFF",X"FFFFFF",X"FEFDF9",X"FFFFFD",X"FBFFFF",X"FAFEFF",X"FDFEFF",X"F4F3F1",X"3D3835",X"070000",X"75051B",X"D80B36",X"CA001F",X"D10624",X"C60021",X"AF102C",X"50081E",X"0F0004",X"362D2E",X"F2E5DD",X"FEFFFA",X"FEFEFF",X"FFFAFF",X"FCFFF6",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFAFF",X"FFF7FF",X"F9FFFF",X"C6C5CB",X"130000",X"543F3C",X"522832",X"321221",X"201011",X"281616",X"2E1221",X"360612",X"000A03",X"301F27",X"000300",X"C7BDBB",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"F9F9F9",X"FDFDFB",X"FFFEFF",X"F6F6EE",X"FFFEFF",X"F2EDEA",X"AFB84F",X"E0E737",X"DDD60C",X"EDE334",X"99A02C",X"060000",X"3D071E",X"871340",X"930020",X"7C070F",X"831828",X"660822",X"F1D3DF",X"F4FDFC",X"FCFEFD",X"F2FEFE",X"F4F9FF",X"F1F7F7",X"FFFEFF",X"FFFDFF",X"FFF9FF",X"D6A8C4",X"35000F",X"4F0022",X"3C0014",X"3B000E",X"4F001F",X"570020",X"5B002E",X"5E0030",X"58002E",X"650041",X"A40561",X"BB0E5E",X"C40962",X"CC0467",X"C51373",X"791055",X"1F001E",X"000D0B",X"001400",X"000F01",X"000E00",X"000E00",X"000B00",X"000E00",X"001505",X"001303",X"000F02",X"001E13",X"001004",X"1BA581",X"36C6A3",X"0C5945",X"040002",X"37153A",X"7B0B6D",X"701179",X"5F0F66",X"41094A",X"2B0F37",X"100C0D",X"070600",X"C5BA3A",X"F9E433",X"DDCB13",X"E0D90D",X"D2D700",X"DCE317",X"C7C429",X"695F06",X"0A0100",X"141011",X"3B4C53",X"312F3D",X"010000",X"8C674A",X"DF8852",X"CE7637",X"D18B67",X"763936",X"000409",X"3B254B",X"9659A9",X"70228F",X"5E047F",X"79118E",X"650078",X"983EAF",X"A63FB2",X"6F0277",X"710075",X"931B97",X"A12BA6",X"75007C",X"710078",X"760078",X"6E0B78",X"82178B",X"801A8A",X"8F2D9C",X"891C99",X"810C90",X"721878",X"300030",X"000102",X"683C21",X"D1692A",X"ED6008",X"F25E00",X"ED6100",X"EC6200",X"F76903",X"F15F09",X"F07225",X"964D1A",X"000100",X"242166",X"4254B6",X"374DA3",X"3A5894",X"090D3C",X"CCD1EE"),
(X"FFF6FE",X"B099A1",X"040000",X"00351F",X"2CCE9C",X"0FD69B",X"00E19C",X"03E9A1",X"00D499",X"08E7A6",X"06E9A2",X"06D994",X"3EDBA4",X"418E7A",X"000012",X"2A0531",X"770574",X"890F96",X"8C0891",X"93029D",X"910985",X"801483",X"3F0B32",X"0D0200",X"1F0100",X"B15B20",X"FF7D15",X"FF7B00",X"FF8A0E",X"F97C0E",X"FA7300",X"FF7C00",X"F7720D",X"FF8E14",X"D6842E",X"5A3C22",X"080004",X"380937",X"6B1070",X"6D017B",X"860E89",X"9C119E",X"8B0B94",X"801599",X"580965",X"1A0027",X"110002",X"833409",X"F38E40",X"E66E0D",X"5A1A00",X"0B0414",X"010002",X"254B72",X"107AE0",X"0075DF",X"097BF7",X"0073E8",X"096ED6",X"1961D0",X"06235F",X"0B0000",X"5C2721",X"CD6F32",X"F97810",X"FA770D",X"F97508",X"F67205",X"F26F03",X"FF8822",X"FB8322",X"EA7518",X"D5641E",X"A44300",X"601400",X"300000",X"200000",X"160000",X"0F0000",X"140B02",X"0F0303",X"150B0A",X"181212",X"171717",X"171D1D",X"182825",X"213832",X"274239",X"242738",X"221C28",X"000208",X"551841",X"BE237F",X"CE0379",X"E40079",X"E60A76",X"DD0185",X"E20082",X"DB087B",X"B3176B",X"57002E",X"190005",X"796F6E",X"FBFFF5",X"FEFEFE",X"F8FAF9",X"FEFFFF",X"FFFFFF",X"FFFAFE",X"FFFEFF",X"FCFFFF",X"F5FFFF",X"DCE4E6",X"386D9F",X"0E71CF",X"0472E3",X"157DEE",X"0064D7",X"0771E7",X"066DE4",X"1170E8",X"0069D9",X"227BE1",X"012B7F",X"545888",X"F1EEF7",X"FFFFF6",X"FAFBF3",X"FCFDFF",X"FFFFFD",X"FFFDF8",X"FFFFFB",X"FDFFFE",X"FAFEFF",X"FDFEFF",X"F3F1F2",X"3A3839",X"000600",X"650F1C",X"CB0F30",X"BE021A",X"CE0C26",X"C30425",X"921527",X"2E0B05",X"0A0000",X"795346",X"FFDFD2",X"FFFFF1",X"F8FFFF",X"FFFBFF",X"FCFFFB",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFB",X"F6F4F7",X"F7FEFF",X"DFC8DC",X"850036",X"C22773",X"C3096C",X"BA0671",X"A60058",X"B21276",X"AA176F",X"691D43",X"000900",X"09204A",X"0072A7",X"A5EBF3",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FDFDFD",X"FFFFFD",X"FFFEFF",X"FFFFF8",X"FFFDFF",X"FFFBFF",X"D9DF95",X"D2D93D",X"E4DE18",X"EAE122",X"CAD248",X"4C4B36",X"340724",X"8A194F",X"96001D",X"9B032C",X"A41E43",X"5C0009",X"C09398",X"FFFEF4",X"FFF8F3",X"FFFEFF",X"FFF8FF",X"F7FFFF",X"FEFCFF",X"FFFDFE",X"F2FFFC",X"EEFAF6",X"7F6A6F",X"290000",X"550715",X"490000",X"43020A",X"3E000A",X"450019",X"390015",X"200111",X"2C0518",X"8A0A3D",X"B5066B",X"CE047E",X"D2007E",X"D00A7B",X"B40B5C",X"7C0034",X"59002A",X"580035",X"5D0029",X"530026",X"50002C",X"540036",X"570034",X"5F0033",X"580032",X"3D0026",X"1B0511",X"0A0406",X"2B8F73",X"29CAA0",X"1CA078",X"001603",X"000012",X"5E2167",X"780387",X"7F0C8F",X"761290",X"4D056B",X"1D002E",X"2D1B1B",X"453F03",X"C5BD5B",X"EAC634",X"D1C32F",X"DCDE61",X"ABAA69",X"1C1210",X"000212",X"001F0E",X"137F45",X"436D7B",X"151531",X"151515",X"A2633A",X"EA6C17",X"E66E00",X"E87822",X"92460A",X"0D0000",X"28021B",X"5C1E5D",X"691877",X"6F087D",X"850687",X"7F0280",X"6C0078",X"70007C",X"7A0184",X"83058A",X"7D0187",X"750084",X"760787",X"861797",X"9B2DAA",X"710083",X"6D0085",X"8819A3",X"9020A6",X"7D008B",X"7C0087",X"6D1272",X"3A0F3C",X"000009",X"250000",X"D16B3A",X"EF6318",X"F9650F",X"EE6109",X"F76B13",X"E45400",X"F46807",X"F27022",X"A0491C",X"060002",X"001054",X"1860C4",X"1166D3",X"1869D5",X"062599",X"B1D5FF"),
(X"FFF9FF",X"AA939B",X"040000",X"3D7862",X"2FD19F",X"0DD499",X"00E5A0",X"00E59D",X"09DDA2",X"05E4A3",X"07EAA3",X"19ECA7",X"30CD96",X"004834",X"000012",X"35103C",X"841281",X"850B92",X"8B0790",X"91009B",X"8E0682",X"770B7A",X"260019",X"0F0402",X"63452B",X"D17B40",X"FF7F17",X"FF8203",X"F78105",X"F77A0C",X"FF7B06",X"FE7800",X"FB7611",X"F98107",X"C5731D",X"180000",X"10030C",X"461745",X"802585",X"7E128C",X"7F0782",X"920794",X"870790",X"7E1397",X"62136F",X"150022",X"160007",X"6D1E00",X"DD782A",X"F27A19",X"591900",X"03000C",X"121013",X"30567D",X"0F79DF",X"0479E3",X"0E80FC",X"1083F8",X"0A6FD7",X"3078E7",X"1A3773",X"0D0000",X"260000",X"BA5C1F",X"FF851D",X"F67309",X"F87407",X"FE7A0D",X"F37004",X"ED6F09",X"E97110",X"F17C1F",X"F5843E",X"E4833F",X"C3773B",X"A56E36",X"8F693C",X"6B5130",X"30210E",X"070000",X"080000",X"080000",X"070101",X"030303",X"000505",X"000A07",X"000F09",X"001007",X"000213",X"100A16",X"000107",X"53163F",X"BC217D",X"D2077D",X"E30078",X"DF036F",X"E5098D",X"E60386",X"D80578",X"B5196D",X"721949",X"310A1D",X"070000",X"C4CABE",X"FFFFFF",X"FBFDFC",X"F9FBFA",X"FFFFFF",X"FFFAFE",X"FEFCFF",X"FBFFFF",X"F7FFFF",X"F9FFFF",X"87BCEE",X"005AB8",X"1583F4",X"066EDF",X"0E77EA",X"046EE4",X"036AE1",X"0C6BE3",X"0771E1",X"0962C8",X"446EC2",X"000434",X"C3C0C9",X"FFFFF6",X"F9FAF2",X"FBFCFF",X"FFFEFC",X"FFFCF7",X"FFFFFB",X"FCFEFD",X"FAFEFF",X"FDFEFF",X"F3F1F2",X"3E3C3D",X"000500",X"6B1522",X"C00425",X"C1051D",X"C6041E",X"C90A2B",X"880B1D",X"210000",X"0E0200",X"946E61",X"FFDFD2",X"FDFFEF",X"F3FDFC",X"FFF9FF",X"FCFFFB",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFA",X"FFFDFF",X"F9FFFF",X"D1BACE",X"8D003E",X"C22773",X"C80E71",X"C7137E",X"BC136E",X"BE1E82",X"B11E76",X"55092F",X"000900",X"2A416B",X"1F97CC",X"9CE2EA",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFFFF",X"FFFFFD",X"FDFCFF",X"FFFFF8",X"FBF9FE",X"FDF8FE",X"FDFFB9",X"D6DD41",X"E0DA14",X"EBE223",X"C7CF45",X"0D0C00",X"5A2D4A",X"AA396F",X"9D0024",X"950026",X"A01A3F",X"790826",X"6B3E43",X"E4DDD3",X"FFFDF8",X"F4F2F5",X"FFF8FF",X"EFFAFC",X"FBF9FC",X"FEFCFD",X"EFFEF9",X"F7FFFF",X"D8C3C8",X"4A0E1A",X"792B39",X"6D1B1F",X"612028",X"5D1229",X"5C1130",X"4D0E29",X"2B0C1C",X"240010",X"800033",X"B90A6F",X"D00680",X"D1007D",X"CC0677",X"BE1566",X"9C1D54",X"7F1D50",X"8A2767",X"882254",X"88255B",X"781E54",X"751D57",X"821F5F",X"871A5B",X"7E2158",X"6E2B57",X"321C28",X"060002",X"268A6E",X"2CCDA3",X"2EB28A",X"1C4D3A",X"2F3044",X"6B2E74",X"7C078B",X"7C098C",X"680482",X"641C82",X"360A47",X"210F0F",X"0E0800",X"554D00",X"F3CF3D",X"E0D23E",X"A5A72A",X"0B0A00",X"0C0200",X"000616",X"367564",X"38A46A",X"47717F",X"070723",X"232323",X"93542B",X"F0721D",X"E36B00",X"E1711B",X"AC6024",X"0A0000",X"1F0012",X"470948",X"6B1A79",X"760F84",X"79007B",X"850886",X"770B83",X"7B0887",X"7C0386",X"7D0084",X"8E1298",X"7E098D",X"720383",X"780989",X"A537B4",X"9923AB",X"75008D",X"72038D",X"6B0081",X"860794",X"A424AF",X"781D7D",X"310633",X"090712",X"2B0000",X"CA6433",X"F3671C",X"F25E08",X"F86B13",X"F1650D",X"F06007",X"EE6201",X"EB691B",X"AE572A",X"201A1C",X"011458",X"145CC0",X"085DCA",X"0C5DC9",X"1534A8",X"B8DCFF"),
(X"F1FFFF",X"959492",X"001805",X"35C190",X"13D99B",X"0BDB9D",X"08E09F",X"00EA9B",X"0BE5AB",X"13D9A8",X"10E1A8",X"3AE1AD",X"39775E",X"000505",X"120427",X"630559",X"9A0698",X"8D058B",X"8F0495",X"8F0C80",X"650C76",X"2E1431",X"0E0000",X"552A00",X"D97D1A",X"F4831D",X"F87A0B",X"FD800A",X"F97B03",X"FF7904",X"FF7A01",X"F97400",X"FF7802",X"F17B0F",X"9D601F",X"0E0200",X"1E001D",X"7B0C73",X"9B0093",X"93008B",X"840391",X"900092",X"8C008E",X"8E0590",X"8E167A",X"310631",X"040004",X"4E1500",X"CB6A25",X"FE8729",X"854716",X"060501",X"020400",X"1F4D71",X"107EE0",X"0576DE",X"0569DB",X"0C82E2",X"1989DD",X"0362DA",X"20528F",X"000A00",X"060200",X"B26D2A",X"F07A10",X"F17708",X"FF810C",X"FD7800",X"F87000",X"FD7100",X"FE7107",X"F86A06",X"F37008",X"FB7A12",X"FC7B15",X"FA7B14",X"FD8622",X"EE8A2C",X"C77624",X"A06114",X"925212",X"803E02",X"621F00",X"460600",X"360000",X"2C0000",X"220000",X"1C0000",X"250000",X"190000",X"000200",X"2A0F1E",X"741D48",X"A91D66",X"CF0A73",X"D20179",X"DF007E",X"DE0385",X"DA0480",X"D60177",X"C91473",X"82174F",X"0F0005",X"7A9285",X"F2F1ED",X"FEFFFD",X"FAFCFB",X"FFFFFF",X"FFFBFF",X"FFFAFE",X"FDFBFC",X"FCFEFB",X"FFFAFF",X"D4E4F3",X"36709E",X"0768C9",X"086FF2",X"1274F3",X"0D77E4",X"0075D2",X"0F73FD",X"006CDB",X"037AD8",X"0875D4",X"003E96",X"425188",X"F2F1FF",X"F9FFFB",X"FBFCFF",X"FEFCFD",X"FFFBF7",X"FFFEF9",X"FDFDFD",X"FCFDFF",X"FEFEFF",X"F3F1F2",X"3D3B48",X"000404",X"6F1129",X"CD002A",X"D30025",X"CC0022",X"C10D34",X"680F21",X"0C0300",X"4B2808",X"C07F57",X"FFE3CE",X"FBFFFA",X"F5FFFF",X"FFFDFD",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFF6F7",X"FEFCFF",X"FCFFFF",X"D9B6CE",X"C60052",X"E21B78",X"DA026D",X"CC026E",X"C6065C",X"CE1177",X"C22389",X"300521",X"0B0109",X"3671B3",X"0099E1",X"B1E0FF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFFFD",X"FDFDFD",X"FCFCFC",X"FFFFF8",X"FBF8FF",X"FCF6FF",X"FFFFDD",X"DDEB93",X"C8CA21",X"EDE427",X"AFAD26",X"0A0800",X"2F1520",X"6A183C",X"88072E",X"9B083E",X"800931",X"5E2F3F",X"070009",X"9A9BB0",X"F6FBFF",X"FFF8FF",X"FCF5ED",X"FFFCFF",X"FFFFFF",X"F4F4F2",X"F8F4F1",X"FFFEFB",X"FDEBE9",X"AC6B73",X"790518",X"A2114A",X"941444",X"A31140",X"A20D37",X"941739",X"5C1E37",X"250E2B",X"691455",X"AF1575",X"C30873",X"C4036C",X"C70867",X"D00561",X"D00E6E",X"C10774",X"D30284",X"C20E69",X"CB076D",X"CB0D7B",X"C61A88",X"C40D81",X"D3037B",X"D00F7C",X"A30863",X"41172B",X"000002",X"217B62",X"25CCA0",X"15B987",X"0A4934",X"392139",X"723674",X"6A027F",X"80038D",X"800591",X"730B84",X"54065C",X"26012A",X"131116",X"060700",X"81755D",X"807A62",X"010800",X"000904",X"003438",X"1D7B7B",X"1C9D8B",X"15AD87",X"248176",X"213239",X"000300",X"A85C2B",X"FF7424",X"E96500",X"FF761C",X"CD6A15",X"2B0000",X"1D030E",X"422251",X"5F0C68",X"800079",X"8B0083",X"7E0084",X"7A098C",X"760684",X"7C0789",X"7A0086",X"840C92",X"7C0B8E",X"861C9A",X"79118C",X"710781",X"7E0E8E",X"790790",X"8B159D",X"7D0183",X"860886",X"901F91",X"651961",X"2A041B",X"1F0000",X"742504",X"DA5E20",X"FF6512",X"FE5D02",X"FF6A0D",X"EF5800",X"FF690F",X"FC6703",X"E86C24",X"A65B3C",X"140A12",X"050239",X"264D9A",X"2660C1",X"286BD4",X"002C98",X"ACE0FF"),
(X"EFFFFD",X"959492",X"0E3926",X"44D09F",X"17DD9F",X"07D799",X"05DD9C",X"00F5A6",X"00DAA0",X"1AE0AF",X"11E2A9",X"22C995",X"00351C",X"000505",X"281A3D",X"76186C",X"950193",X"8E068C",X"900596",X"931084",X"5A016B",X"150018",X"100000",X"855A25",X"E68A27",X"EB7A14",X"F17304",X"F67903",X"FD7F07",X"FF7803",X"FC7100",X"FB7600",X"FF7600",X"F17B0F",X"7F4201",X"0A0000",X"2C0A2B",X"7A0B72",X"9D0095",X"95008D",X"81008E",X"950097",X"950797",X"900792",X"830B6F",X"3F143F",X"040004",X"511800",X"D77631",X"F98224",X"995B2A",X"010000",X"090B06",X"0A385C",X"0C7ADC",X"097AE2",X"1074E6",X"0074D4",X"0A7ACE",X"0F6EE6",X"154784",X"011305",X"040000",X"AE6926",X"F88218",X"EE7405",X"FB7C07",X"FA7500",X"FD7500",X"FE7201",X"FF7309",X"F96B07",X"F9760E",X"FF7E16",X"FE7D17",X"F67710",X"EF7814",X"E37F21",X"D58432",X"CA8B3E",X"CE8E4E",X"C9874B",X"C17E49",X"BB7B4F",X"B57954",X"A2704F",X"815838",X"654222",X"51271B",X"230200",X"040601",X"110005",X"49001D",X"9D115A",X"D00B74",X"D90880",X"E80087",X"E4098B",X"D7017D",X"E10C82",X"C40F6E",X"90255D",X"321A28",X"000900",X"D1D0CC",X"FEFFFD",X"FBFDFC",X"FBFBFD",X"FFFDFF",X"FFFDFF",X"FFFDFE",X"FAFCF9",X"FFF5FD",X"F2FFFF",X"77B1DF",X"0465C6",X"0C73F6",X"0E70EF",X"036DDA",X"0076D3",X"096DF7",X"0571E0",X"0071CF",X"0370CF",X"2969C1",X"000D44",X"B1B0BE",X"F8FFFA",X"FBFCFF",X"FEFCFD",X"FFFAF6",X"FFFEF9",X"FDFDFD",X"FCFDFF",X"FEFEFF",X"F3F1F2",X"393744",X"000404",X"6A0C24",X"D60433",X"D30025",X"D10027",X"BD0930",X"650C1E",X"070000",X"735030",X"CB8A62",X"FFDFCA",X"F9FFF8",X"F7FFFF",X"FFFDFD",X"FCFCFC",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFCFD",X"FDFBFE",X"F7FAFF",X"DAB7CF",X"CC0258",X"E01976",X"DA026D",X"CF0571",X"CB0B61",X"C5086E",X"A90A70",X"29001A",X"070005",X"4B86C8",X"02A3EB",X"ABDAFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FDFCFF",X"FFFFFD",X"FDFDFD",X"FFFFFF",X"FFFFF8",X"FFFDFF",X"FFFCFF",X"FFFFDB",X"F6FFAC",X"D9DB32",X"EAE124",X"C8C63F",X"2E2C13",X"110002",X"5F0D31",X"8E0D34",X"910034",X"760027",X"1F0000",X"140816",X"020318",X"E4E9FC",X"FFF1FD",X"FFFEF6",X"FBF4FC",X"FEFEFF",X"FAFAF8",X"FFFEFB",X"FBF7F4",X"FFFAF8",X"FFC0C8",X"750114",X"9D0C45",X"8A0A3A",X"9E0C3B",X"99042E",X"8F1234",X"571932",X"17001D",X"580344",X"B31979",X"C70C77",X"D11079",X"D11271",X"CB005C",X"D10F6F",X"C60C79",X"D10082",X"BC0863",X"D20E74",X"BF016F",X"AE0270",X"BD067A",X"CA0072",X"C2016E",X"A80D68",X"42182C",X"010103",X"1B755C",X"20C79B",X"12B684",X"003924",X"0E000E",X"350037",X"740C89",X"850892",X"79008A",X"6E067F",X"66186E",X"310C35",X"030106",X"101109",X"0B0000",X"0D0700",X"121907",X"132E29",X"2E686C",X"45A3A3",X"22A391",X"039B75",X"217E73",X"102128",X"070A00",X"9D5120",X"FD7020",X"E96500",X"F4670D",X"D97621",X"754541",X"110002",X"1C002B",X"5B0864",X"84007D",X"8C0084",X"810287",X"7C0B8E",X"891997",X"7A0587",X"7B0187",X"8B1399",X"720184",X"67007B",X"69017C",X"6E047E",X"790989",X"78068F",X"901AA2",X"85098B",X"7E007E",X"7D0C7E",X"60145C",X"220013",X"350B00",X"A25332",X"F27638",X"FD620F",X"FF670C",X"F45900",X"FC650A",X"FB6107",X"FA6501",X"EB6F27",X"AB6041",X"090007",X"09063D",X"2B529F",X"2761C2",X"1B5EC7",X"0E3DA9",X"ABDFFF"),
(X"FCFFFD",X"928A88",X"05945F",X"2AD89D",X"06D293",X"1AD59E",X"0DE2A0",X"03E59D",X"00E592",X"0AD691",X"4CE4B5",X"2F8268",X"000404",X"290426",X"5F0E5D",X"8B0F87",X"9100A5",X"9701A0",X"920B81",X"6E0D76",X"270221",X"190200",X"793E00",X"E57424",X"FF7301",X"FE7B0F",X"F1710E",X"F8690B",X"FF7110",X"FD6F09",X"F36D0A",X"FF7A1E",X"F9710D",X"E8741D",X"87461C",X"0D0000",X"27042E",X"731273",X"88098E",X"7C0A84",X"860691",X"920093",X"980496",X"960795",X"91137E",X"380A3B",X"07000B",X"622103",X"D27629",X"FF8E26",X"C75810",X"1B0000",X"1F1122",X"010012",X"37577E",X"3A76B2",X"3165BB",X"2E70D0",X"3A78CD",X"3366C2",X"131B42",X"250C07",X"200000",X"CE6514",X"FF7A07",X"FF7903",X"FF7A00",X"F66F00",X"F67000",X"FF800C",X"FA7A0D",X"F77811",X"F67E03",X"F17E0B",X"ED7C12",X"F17B17",X"F77912",X"FE7608",X"FF7300",X"FF7200",X"FA7E02",X"FE7D06",X"FF7A0E",X"FF7713",X"FC751B",X"F87821",X"F27A24",X"ED7924",X"C17F35",X"66300A",X"0B0000",X"120A15",X"0B0004",X"4A0E27",X"AC1C62",X"BE0D75",X"F7037F",X"EE0280",X"E1007D",X"DE027E",X"DC077B",X"BF106D",X"6C0E43",X"0D000C",X"827D7A",X"F9F8F6",X"FBFDFC",X"FFFFFF",X"FFFAFE",X"FDF7F9",X"FFFEFB",X"FBFAF5",X"FDF4FF",X"FFFEFF",X"D7EAF1",X"1C5688",X"297DE0",X"0968E0",X"026DE1",X"0078E2",X"076BE3",X"076BE3",X"0877E2",X"0175D8",X"0F69D9",X"0F3AAD",X"41539B",X"DCF2FF",X"FBFFFF",X"FBFBFD",X"FFFEFB",X"FAF6F3",X"FFFFFD",X"FEFFFF",X"F8F8FA",X"F6F4F5",X"473040",X"030305",X"630A1C",X"C4042B",X"CD0625",X"C30423",X"AE0F2F",X"520815",X"030007",X"B1633C",X"D1803E",X"FEEBCB",X"F5FFFF",X"F8FDFF",X"FFFFF5",X"FFFCFD",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"F7FFFA",X"FFFEFB",X"FFF5FF",X"E79FC5",X"D90064",X"DB1C84",X"D6027A",X"D10078",X"DC0876",X"C5127A",X"680E42",X"00000B",X"092145",X"269EDB",X"00A4E0",X"B7D6FF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFFFB",X"FFFEFF",X"FEFFFD",X"FFFFF8",X"FEFDFF",X"FFFCFF",X"FFFEF2",X"F8FFF1",X"E8EB84",X"DFD849",X"CBC54B",X"352F0D",X"250D0B",X"782D4B",X"84082C",X"761828",X"400815",X"000315",X"07316B",X"002E8A",X"77A8F5",X"EBFFFF",X"E8FFE7",X"FFF6FD",X"FEFDFB",X"FAFFF9",X"FCFBF9",X"FFFEFF",X"FCF8F7",X"FFEAED",X"B88187",X"730522",X"83203D",X"8B1F41",X"831B3C",X"7E1E39",X"5A222D",X"010000",X"2D161E",X"693355",X"75284A",X"762A46",X"772848",X"862254",X"8A275E",X"8E3062",X"931F50",X"A51C60",X"C90C68",X"D90372",X"C80175",X"C20073",X"D70479",X"CE0B74",X"AA0D64",X"591136",X"160410",X"12644E",X"25C79E",X"2EB896",X"0F4839",X"02000E",X"1A1035",X"6D0C73",X"850784",X"931799",X"780D81",X"62035D",X"3B043B",X"0A0015",X"1C0521",X"021911",X"010E14",X"3F5664",X"347F84",X"109E8E",X"009D83",X"1BB4A2",X"1F9795",X"12795C",X"030400",X"331800",X"BC5E2A",X"FC711E",X"F7720B",X"F75807",X"F8752F",X"C6662C",X"240000",X"100604",X"240A39",X"611F76",X"6F1078",X"770C74",X"79066E",X"6C0973",X"89228F",X"87198A",X"811084",X"6F0275",X"A53EAB",X"9F35A1",X"730870",X"8A007E",X"8E048B",X"880788",X"750374",X"6B1472",X"4E125C",X"320732",X"1A0000",X"6A2100",X"D87635",X"E05F0B",X"FD6B08",X"F56200",X"F16300",X"F06805",X"F76C0D",X"E95E00",X"FF7331",X"AC5037",X"000203",X"0F1340",X"263379",X"354E9E",X"326AB7",X"0D3479",X"BDE4FF"),
(X"FAFFFB",X"A29A98",X"19A873",X"32E0A5",X"09D596",X"1AD59E",X"0ADF9D",X"00E29A",X"00DF8C",X"24F0AB",X"38D0A1",X"00442A",X"000505",X"421D3F",X"671665",X"870B83",X"8D00A1",X"9903A2",X"960F85",X"5B0063",X"170011",X"1F0800",X"BB803C",X"F48333",X"FF7301",X"FB780C",X"F2720F",X"FB6C0E",X"FF7110",X"FF710B",X"F16B08",X"F36C10",X"FF7713",X"F5812A",X"9D5C32",X"0D0000",X"200027",X"6B0A6B",X"8B0C91",X"82108A",X"870792",X"980099",X"960294",X"90018F",X"860873",X"360839",X"0A000E",X"6F2E10",X"DC8033",X"FF8018",X"E6772F",X"472219",X"0B000E",X"040015",X"000930",X"003B77",X"164AA0",X"185ABA",X"1A58AD",X"093C98",X"00072E",X"120000",X"4E2020",X"DD7423",X"FE7704",X"F87000",X"FF7800",X"FF7F02",X"FF830A",X"FF7D09",X"FA7A0D",X"FF8019",X"FB8308",X"F78411",X"F38218",X"F27C18",X"F2740D",X"F87002",X"FF7300",X"FF7801",X"F47800",X"F77600",X"FA7307",X"F9710D",X"F77016",X"F1711A",X"EB731D",X"E8741F",X"D9974D",X"97613B",X"0A0000",X"160E19",X"1F0E18",X"280005",X"8D0043",X"C8177F",X"ED0075",X"EA007C",X"E3017F",X"E10581",X"DA0579",X"BC0D6A",X"76184D",X"230D22",X"040000",X"DAD9D7",X"FAFCFB",X"FAFAFC",X"FFFAFE",X"FFFDFF",X"FFFDFA",X"FFFEF9",X"FFF9FF",X"FFFEFF",X"E8FBFF",X"79B3E5",X"0051B4",X"207FF7",X"0D78EC",X"0076E0",X"076BE3",X"0B6FE7",X"0372DD",X"006BCE",X"0B65D5",X"4873E6",X"001159",X"AAC0CE",X"F8FDFF",X"F8F8FA",X"FFFEFB",X"FFFDFA",X"F6F6F4",X"FCFDFF",X"FFFFFF",X"EFEDEE",X"493242",X"000002",X"630A1C",X"C8082F",X"CD0625",X"C90A29",X"B01131",X"47000A",X"0A040E",X"C3754E",X"DE8D4B",X"FCE9C9",X"EFFCFF",X"F6FBFE",X"FFFFF6",X"FFF9FA",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"F3FFF6",X"FEFAF7",X"FFF6FF",X"EAA2C8",X"D50060",X"D81981",X"D6027A",X"D90480",X"D5016F",X"C7147C",X"6B1145",X"01000C",X"2B4367",X"33ABE8",X"00A6E2",X"B6D5FF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFFFB",X"FFFEFF",X"FEFFFD",X"FFFFF8",X"FEFDFF",X"FFFCFF",X"FFFEF2",X"F7FFF0",X"FDFF99",X"EDE657",X"C9C349",X"0F0900",X"2E1614",X"671C3A",X"8B0F33",X"731525",X"3B0310",X"041527",X"1A447E",X"3362BE",X"2B5CA9",X"C3DBF7",X"F0FFEF",X"FFF8FF",X"FCFBF9",X"FCFFFB",X"FEFDFB",X"FAF8F9",X"FDF9F8",X"FFF7FA",X"FFCBD1",X"730522",X"670421",X"7F1335",X"700829",X"5F001A",X"330006",X"272622",X"0F0000",X"22000E",X"4C0021",X"420012",X"3E000F",X"5B0029",X"66033A",X"57002B",X"7A0637",X"84003F",X"BF025E",X"D6006F",X"C50072",X"C70578",X"D50277",X"C5026B",X"AA0D64",X"60183D",X"180612",X"055741",X"23C59C",X"34BE9C",X"366F60",X"00000C",X"271D42",X"74137A",X"830582",X"84088A",X"7E1387",X"72136D",X"440D44",X"22122D",X"3A233F",X"000901",X"000309",X"253C4A",X"358085",X"20AE9E",X"00AB91",X"0EA795",X"39B1AF",X"1D8467",X"020300",X"5F4429",X"C46632",X"FF7926",X"EF6A03",X"FF600F",X"E96620",X"DA7A40",X"64370D",X"0B0100",X"19002E",X"55136A",X"771880",X"80157D",X"7E0B73",X"68056F",X"8C2592",X"942697",X"750478",X"75087B",X"A13AA7",X"A238A4",X"6D026A",X"89007D",X"90068D",X"7A007A",X"861485",X"6C1573",X"3C004A",X"240024",X"310E15",X"A9602D",X"DD7B3A",X"E86713",X"EC5A00",X"FF6F07",X"F46600",X"EF6704",X"EC6102",X"FD7209",X"ED5F1D",X"953920",X"616566",X"373B68",X"000046",X"0E2777",X"0F4794",X"062D72",X"B6DDFE"),
(X"FBFAF8",X"8EB7A5",X"00C779",X"0DE39B",X"0CCF93",X"07E2A0",X"06E69F",X"15E29D",X"25E59C",X"41C395",X"30655B",X"000013",X"30083C",X"770D6F",X"910089",X"9404A1",X"870492",X"840C78",X"5D1561",X"21111E",X"190000",X"9C3C00",X"FF8933",X"F38C15",X"EC9039",X"D48A31",X"E2994A",X"F39A58",X"E1823E",X"E5872F",X"FC8C20",X"FF7200",X"F4690C",X"F87A14",X"BC672E",X"160000",X"15031D",X"4F1349",X"820F76",X"8A0085",X"80088E",X"940099",X"900296",X"841099",X"61176E",X"1B0D26",X"0C0000",X"863E03",X"F29420",X"F37D02",X"FE8C19",X"AF621A",X"270000",X"3E0E0C",X"391517",X"0D0010",X"0C0000",X"040000",X"070000",X"0D0000",X"2B0000",X"561000",X"B85D28",X"FC821D",X"FF7512",X"FD7813",X"FA7C18",X"ED7B1A",X"EE8B2D",X"E28D33",X"DD923F",X"CB8638",X"9F6744",X"B07145",X"C87D3C",X"E0822B",X"F17F1C",X"FA7B14",X"F97513",X"F47117",X"FC770E",X"FC740E",X"FF720E",X"FF7312",X"FF7212",X"FF710D",X"FC730B",X"FD760D",X"EF8B2B",X"8D4714",X"070400",X"265359",X"045747",X"001300",X"390E21",X"76204F",X"AF1D66",X"D30D6E",X"DF0172",X"D30979",X"D60A79",X"DF0774",X"BA1066",X"731248",X"110303",X"7A7172",X"FBF9FA",X"FBFBFB",X"FFFEFF",X"FFFBFD",X"FAF4F4",X"FFFBF8",X"FCF6FA",X"F7F5F8",X"FFFFFD",X"DEECED",X"315F80",X"1E70C2",X"1B78EF",X"1265E9",X"0D73E2",X"016BDB",X"0F72E7",X"0F62E2",X"1263E8",X"1B6EE8",X"165ABD",X"2A58A6",X"E9F3FD",X"FBFFFF",X"F6F4F5",X"FFFDFA",X"FCFCFC",X"FEFEFF",X"FFFFFF",X"EBE9EA",X"483E3C",X"040000",X"5E1318",X"B6172D",X"B90C1F",X"B11B27",X"851D24",X"220000",X"400600",X"F06D27",X"EF8726",X"FFEBB6",X"FAF8FD",X"FFFDFE",X"FBFFF8",X"FDF8FF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FBFFFB",X"F8FAF5",X"FFF6F9",X"EE9CC2",X"C7005A",X"D0217E",X"C30A6F",X"C10D70",X"D7096E",X"A11C6B",X"282104",X"000309",X"1579AB",X"1FB7E8",X"009CD5",X"AFDFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFFFA",X"FFFEFF",X"FEFFFD",X"FEFFFA",X"FEFDFF",X"FEFEFE",X"FEFBFF",X"FFFBFF",X"FBFADB",X"E1E19B",X"C9CA6C",X"463E1A",X"190000",X"671138",X"8D0722",X"550F19",X"0F0000",X"1E223D",X"2F5EA2",X"2367D2",X"1453BC",X"6EA7DE",X"EAFDFF",X"F8FEFC",X"F5F4F0",X"FAFCF7",X"F5FFFF",X"F5FFFF",X"FFFBFF",X"FFFDFF",X"F5FBF7",X"B48A94",X"120000",X"25130F",X"040400",X"170400",X"2A0B00",X"3F3800",X"543700",X"0F0300",X"150000",X"1B0400",X"0F0000",X"190900",X"0D0100",X"110500",X"160012",X"1E001B",X"851152",X"C40A6D",X"C90372",X"D30E81",X"D3077A",X"C10069",X"B7126E",X"6B1D47",X"000105",X"17624E",X"22C49D",X"18CC9D",X"0B7A59",X"00030A",X"3C3E57",X"662583",X"6D0077",X"7B028D",X"750188",X"7A0379",X"530A53",X"19021F",X"36192B",X"641A2B",X"38050E",X"060000",X"134539",X"29937D",X"15A58A",X"0AAA92",X"12B69E",X"0A8B65",X"001319",X"110002",X"86442C",X"DF772E",X"EA7504",X"FB6300",X"FF6D06",X"FF6411",X"E56422",X"611200",X"160000",X"190A0F",X"381237",X"551854",X"622068",X"7A168A",X"7F138D",X"800B8D",X"8E169B",X"7B0388",X"750082",X"720079",X"820A86",X"67207E",X"531373",X"5D2677",X"421745",X"2B1023",X"260E0C",X"240000",X"84370B",X"ED7624",X"EF6C14",X"FD6A0A",X"EE5500",X"FF7309",X"F56800",X"F16300",X"F36503",X"F5690A",X"E4753D",X"622415",X"5C5354",X"53293D",X"16000A",X"230F32",X"1D204D",X"000215",X"C4D2DF"),
(X"FFFFFD",X"A0C9B7",X"00D385",X"0EE49C",X"1ADDA1",X"13EEAC",X"08E8A1",X"15E29D",X"2DEDA4",X"159769",X"001107",X"222538",X"50285C",X"841A7C",X"A4109C",X"A111AE",X"9C19A7",X"951D89",X"4B034F",X"1F0F1C",X"35120C",X"D27236",X"FF8630",X"F79019",X"DB7F28",X"B66C13",X"A35A0B",X"B75E1C",X"D37430",X"E78931",X"F7871B",X"FF7B03",X"F86D10",X"FC7E18",X"D07B42",X"29090C",X"1F0D27",X"50144A",X"8E1B82",X"9E1299",X"8E169C",X"A30EA8",X"9E10A4",X"9723AC",X"641A71",X"1B0D26",X"23160E",X"BD753A",X"E28410",X"FF9116",X"F3810E",X"D98C44",X"9D6856",X"643432",X"351113",X"0D0010",X"231709",X"1B170B",X"181101",X"210E10",X"5D3011",X"BA7436",X"E48954",X"F07611",X"FF7613",X"FF821D",X"FF8622",X"F38120",X"F79436",X"DB862C",X"BB701D",X"803B00",X"3E0600",X"4B0C00",X"7F3400",X"CC6E17",X"FC8A27",X"FE7F18",X"F77311",X"F9761C",X"FE7910",X"FB730D",X"FF710D",X"FF7514",X"FF7414",X"FF720E",X"FD740C",X"FF7910",X"E27E1E",X"7C3603",X"050200",X"346167",X"55A898",X"1D543F",X"200008",X"5E0837",X"B3216A",X"E01A7B",X"F01283",X"E01686",X"E01483",X"EA127F",X"C71D73",X"86255B",X"302222",X"0E0506",X"D6D4D5",X"FDFDFD",X"FDF9FA",X"FBF5F7",X"FFFDFD",X"FFFBF8",X"FDF7FB",X"FFFDFF",X"F8F8F6",X"F0FEFF",X"90BEDF",X"004EA0",X"217EF5",X"186BEF",X"1076E5",X"0973E3",X"187BF0",X"176AEA",X"1768ED",X"1E71EB",X"3579DC",X"154391",X"9EA8B2",X"FBFFFF",X"FDFBFC",X"F8F4F1",X"FDFDFD",X"FBFBFD",X"FCFCFE",X"F7F5F6",X"443A38",X"0A0600",X"6A1F24",X"BE1F35",X"C4172A",X"B8222E",X"80181F",X"220000",X"814733",X"FF7E38",X"EB8322",X"FFECB7",X"FFFDFF",X"FCFAFB",X"FBFFF8",X"FFFDFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FBFFFB",X"FAFCF7",X"FFF6F9",X"ED9BC1",X"CC035F",X"D82986",X"CE157A",X"CB177A",X"E11378",X"95105F",X"1F1800",X"101D23",X"399DCF",X"20B8E9",X"0096CF",X"ABDBFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFFFA",X"FFFEFF",X"FEFFFD",X"FEFFFA",X"FEFDFF",X"FEFEFE",X"FEFBFF",X"F9F2FF",X"FFFFE3",X"FFFFBF",X"D0D173",X"352D09",X"48282D",X"8A345B",X"A01A35",X"5B151F",X"2B1517",X"040823",X"2E5DA1",X"2D71DC",X"2362CB",X"276097",X"CFE2F3",X"FBFFFF",X"FFFFFB",X"F7F9F4",X"F4FFFE",X"F5FFFF",X"FFFCFF",X"FFF9FD",X"FBFFFD",X"FFD8E2",X"5C4245",X"362420",X"44442A",X"8D7A52",X"B3945B",X"A8A151",X"B19446",X"ADA167",X"AD966D",X"8E7757",X"908158",X"847443",X"776B41",X"4C4034",X"22091E",X"250222",X"871354",X"C3096C",X"C1006A",X"C40072",X"C8006F",X"C00068",X"BB1672",X"63153F",X"000408",X"196450",X"29CBA4",X"0BBF90",X"2B9A79",X"00070E",X"000018",X"4E0D6B",X"7E0F88",X"860D98",X"841097",X"7D067C",X"4B024B",X"2B1431",X"371A2C",X"722839",X"35020B",X"100806",X"001004",X"157F69",X"22B297",X"07A78F",X"00A088",X"21A27C",X"12252B",X"0F0000",X"5F1D05",X"D97128",X"E26D00",X"FF6B00",X"F66300",X"F15603",X"F1702E",X"B5663B",X"2C1000",X"0A0000",X"220021",X"2F002E",X"3A0040",X"600070",X"851993",X"881395",X"870F94",X"740081",X"830E90",X"7C0583",X"7F0783",X"5D1674",X"551575",X"450E5F",X"28002B",X"110009",X"160000",X"9B6D55",X"C27549",X"E06917",X"E25F07",X"F66303",X"F96000",X"FE6A00",X"F66900",X"EF6100",X"F76907",X"F06405",X"D1622A",X"4D0F00",X"060000",X"481E32",X"331227",X"321E41",X"212451",X"000A1D",X"C6D4E1"),
(X"EBFFFF",X"8FD9BE",X"1BC086",X"1BC98E",X"30C196",X"1ED39C",X"1FC891",X"2EC892",X"299677",X"000106",X"08000D",X"07011D",X"64105B",X"760C6E",X"5E0C70",X"780A7A",X"5F0D57",X"4E1245",X"060002",X"000A00",X"694C22",X"D87645",X"E78B3E",X"A17826",X"070506",X"030000",X"030004",X"04020F",X"01000C",X"332117",X"986236",X"E58E47",X"E26B17",X"DA720F",X"B86C30",X"250400",X"030000",X"130014",X"530A59",X"780982",X"700D6A",X"7F0A75",X"7A0669",X"6A106A",X"30002C",X"110000",X"3B0E08",X"CB7B3E",X"E77B23",X"D87321",X"DA7A13",X"E2830F",X"E3852E",X"B96E2A",X"AA661F",X"A65617",X"BE6D3E",X"A75617",X"A1520F",X"BC6635",X"CB7834",X"E08723",X"E06E0E",X"E58018",X"DA7C1C",X"D0781F",X"C47731",X"A06432",X"673E22",X"120000",X"060000",X"01010B",X"070002",X"060007",X"070007",X"150000",X"592913",X"AF6631",X"DA7F2C",X"DA7614",X"E47524",X"E17020",X"E37020",X"E87323",X"E87421",X"E37119",X"E37216",X"E67819",X"D8834D",X"6F3E1E",X"000400",X"0B3E3F",X"4AAB98",X"298266",X"000500",X"000002",X"4B0424",X"950F4A",X"C11061",X"BF0E66",X"B80A63",X"BD045F",X"B60B5A",X"960E4E",X"220D12",X"0A0000",X"736F6E",X"F4F3F1",X"FFFFFD",X"FDF9FA",X"FFFDFF",X"FAF8FB",X"FFFFF7",X"FEFFFF",X"FFFBFF",X"FFFEF8",X"E7F3F3",X"4C7595",X"174C90",X"2B59B1",X"0E5FB8",X"075DA6",X"105DAD",X"1857C0",X"1558C0",X"1366B4",X"05559C",X"1753AB",X"203040",X"D5DDE8",X"FEFFFF",X"F9F7F8",X"FCFCFC",X"FAFAFC",X"FBF9FC",X"FBF7F8",X"09140C",X"060000",X"4C0813",X"910721",X"A00620",X"81111D",X"350906",X"000200",X"A15D36",X"E27A3B",X"CD7F34",X"FCE6B7",X"FFFDF8",X"FCFAFB",X"F6FFFA",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFF8FF",X"F3FFFF",X"F2FBFF",X"DF93BA",X"AB0655",X"B81669",X"B30A5B",X"B41059",X"8B114A",X"39012E",X"000600",X"010B40",X"1376C7",X"1B8ECD",X"178DBD",X"9DE5FD",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFD",X"FFFFF8",X"FFFDFF",X"FEFFFD",X"FEFFFB",X"FDFEFF",X"FEFFF7",X"FDFBFF",X"FFFAFF",X"F6F8F3",X"EFF5E7",X"DFE0B6",X"0D0300",X"0D0000",X"37031A",X"58020F",X"460D20",X"100004",X"07000B",X"071230",X"153463",X"2A4D83",X"00214B",X"77729B",X"E7F1F0",X"FFFFFD",X"FEFAF9",X"FCFFFF",X"FBFCFF",X"FFF6FF",X"FFF9FF",X"FEFFFF",X"FFFFF8",X"D2CEB1",X"9D8D4F",X"B7AE45",X"D8B93C",X"C9A11E",X"B7A622",X"D3A837",X"D0B00D",X"D1B428",X"CEA730",X"DBB634",X"CCB823",X"D2C042",X"B99F64",X"371D1C",X"1D202F",X"712A56",X"B82B77",X"C6267E",X"C62380",X"CF2182",X"D22483",X"CC2984",X"922054",X"200F19",X"31554B",X"2DB795",X"10D7A0",X"20C18D",X"304945",X"332C3E",X"493477",X"6B207D",X"7B2890",X"74218B",X"87258A",X"6F3776",X"2D293A",X"322225",X"A2203C",X"893042",X"431A22",X"261D20",X"212C30",X"4D827A",X"289B7E",X"18BE8E",X"16A683",X"144E52",X"182939",X"130E0B",X"A87351",X"E78846",X"E66A12",X"EC6C09",X"F67C26",X"F46C20",X"F06B26",X"D56F2D",X"8D4811",X"2B0000",X"371E17",X"2A282D",X"2E2135",X"402C47",X"4D3255",X"4F3059",X"5D4169",X"553B60",X"4D3253",X"492C4B",X"35263B",X"281F34",X"2A1921",X"200000",X"723310",X"A04F22",X"F17C46",X"FF7632",X"EB6A19",X"EA6614",X"EB6412",X"F5711E",X"F0721D",X"F1751F",X"EE6D1A",X"ED6917",X"EC7D4F",X"795535",X"111610",X"402B32",X"951F2F",X"A53436",X"7A202A",X"893E5D",X"060000",X"D6D0D0"),
(X"E5FFF9",X"A1EBD0",X"3EE3A9",X"3AE8AD",X"4CDDB2",X"38EDB6",X"3FE8B1",X"55EFB9",X"3EAB8C",X"66696E",X"68606D",X"7A7490",X"A7539E",X"BF55B7",X"AB59BD",X"BF51C1",X"AC5AA4",X"93578A",X"6D6469",X"5D6A60",X"B6996F",X"FB9968",X"F29649",X"9F7624",X"666465",X"7C7877",X"7C777D",X"72707D",X"6E6C79",X"6F5D53",X"986236",X"DE8740",X"FF9844",X"FF9835",X"E4985C",X"86655C",X"6B6768",X"735D74",X"9E55A4",X"B647C0",X"B754B1",X"C651BC",X"C04CAF",X"AF55AF",X"895885",X"785F65",X"946761",X"EB9B5E",X"FD9139",X"FF9A48",X"FFA63F",X"FB9C28",X"F99B44",X"F0A561",X"EFAB64",X"EC9C5D",X"E29162",X"F1A061",X"EE9F5C",X"EC9665",X"ED9A56",X"F19834",X"FF8E2E",X"F9942C",X"F79939",X"F69E45",X"D88B45",X"9A5E2C",X"7C5337",X"705A4F",X"756C6F",X"63636D",X"71666C",X"716772",X"716571",X"765C5D",X"885842",X"AE6530",X"E08532",X"FFA240",X"FD8E3D",X"FC8B3B",X"FE8B3B",X"FF8D3D",X"FF8E3B",X"FF8D35",X"FF8E32",X"FF9132",X"EA955F",X"9D6C4C",X"57625A",X"588B8C",X"58B9A6",X"67C0A4",X"83928B",X"656567",X"914A6A",X"D6508B",X"FD4C9D",X"FA49A1",X"F84AA3",X"FF48A3",X"FD52A1",X"E25A9A",X"867176",X"7E6F72",X"858180",X"EFEEEC",X"FFFFFD",X"FFFBFC",X"FCF7FB",X"F9F7FA",X"FCFCF4",X"F9FAFE",X"FFFDFF",X"FFFBF5",X"F4FFFF",X"ABD4F4",X"487DC1",X"6492EA",X"4899F2",X"4399E2",X"4794E4",X"5291FA",X"5497FF",X"4194E2",X"4898DF",X"5793EB",X"566676",X"CCD4DF",X"FAFBFF",X"FFFDFE",X"FFFFFF",X"FCFCFE",X"FCFAFD",X"F6F2F3",X"667169",X"6D6562",X"A35F6A",X"D94F69",X"EA506A",X"CC5C68",X"8D615E",X"696C61",X"CA865F",X"FC9455",X"EFA156",X"FFEBBC",X"FFFDF8",X"FEFCFD",X"F8FFFC",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFF8FF",X"F4FFFF",X"F2FBFF",X"F4A8CF",X"E64190",X"EC4A9D",X"EE4596",X"EB4790",X"D25891",X"98608D",X"60716B",X"757FB4",X"50B3FF",X"48BBFA",X"3EB4E4",X"96DEF6",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFD",X"FFFFF8",X"FFFDFF",X"FEFFFD",X"FEFFFB",X"FDFEFF",X"FEFFF7",X"FDFBFF",X"FFF7FF",X"FEFFFB",X"F9FFF1",X"FBFCD2",X"948A80",X"715E60",X"9B677E",X"B15B68",X"A2697C",X"7E6972",X"716475",X"5C6785",X"436291",X"4C6FA5",X"5679A3",X"524D76",X"D3DDDC",X"FCFBF9",X"FCF8F7",X"FCFFFF",X"FDFEFF",X"FFF8FF",X"FFF9FF",X"F9FBFA",X"FCFCF4",X"FDF9DC",X"E1D193",X"B6AD44",X"C5A629",X"DDB532",X"BDAC28",X"CA9F2E",X"D9B916",X"AE9105",X"C09922",X"BC9715",X"C4B01B",X"B8A628",X"C1A76C",X"1D0302",X"00000E",X"400025",X"8D004C",X"A6065E",X"A4015E",X"AE0061",X"B00261",X"9F0057",X"700032",X"0D0006",X"000F05",X"1AA482",X"00C28B",X"01A26E",X"000804",X"03000E",X"140042",X"4B005D",X"4C0061",X"500067",X"540057",X"25002C",X"040011",X"0C0000",X"760010",X"6A1123",X"200000",X"060000",X"000307",X"001810",X"0F8265",X"009D6D",X"0A9A77",X"053F43",X"000313",X"040000",X"380300",X"B45513",X"D55901",X"E06000",X"D25802",X"E45C10",X"DF5A15",X"B95311",X"B9743D",X"815332",X"150000",X"010004",X"07000E",X"0B0012",X"0F0017",X"15001F",X"1C0028",X"150020",X"0F0015",X"110013",X"08000E",X"0C0318",X"120109",X"320800",X"A46542",X"C37245",X"BD4812",X"E54C08",X"DA5908",X"DB5705",X"D95200",X"DB5704",X"D85A05",X"D45802",X"DE5D0A",X"D85402",X"992A00",X"230000",X"000200",X"1C070E",X"7C0616",X"680000",X"5D030D",X"590E2D",X"110A02",X"D5CFCF"),
(X"FDFFFE",X"FFF6F8",X"EEF7F2",X"FEF9FD",X"E4FFFE",X"FCF7FE",X"E5F8F2",X"E8FCF1",X"EEFAF8",X"F6F9F2",X"FFF4EF",X"FFF4FA",X"FFECFF",X"FFEAFF",X"F9EDF7",X"F5FAF3",X"FAEDFF",X"FBEDFA",X"FFF8FF",X"FCEFF6",X"F4EDE3",X"FFFFDC",X"FAF2DF",X"FFEFFA",X"F6FAFF",X"FFF1FC",X"FFF0FC",X"FCF9FF",X"F5F9FF",X"FBF3FF",X"FFF3F4",X"FFF7E9",X"FAF1E8",X"F9EFE3",X"FFF0F3",X"FEEFF6",X"FFFDEE",X"FAFDF2",X"FBF9FF",X"F8ECF8",X"F4F1FA",X"F9EEFE",X"FAEDF6",X"FAF2FF",X"F5F9FC",X"FDF7FF",X"FDE6FF",X"FFEFDB",X"F5F3E6",X"FDF2EC",X"F2F4E7",X"F4FAF0",X"FFF0F2",X"FAE6DF",X"F7F4E1",X"F9F9F1",X"EFF0E2",X"FFF0F0",X"FEF0EF",X"FFEFE1",X"F7F5E6",X"F4E8E8",X"FFE8EC",X"F2FAEB",X"FFF4E0",X"F9EDDD",X"FBF1E8",X"FDF1F1",X"FFF5F9",X"FEF5FA",X"FBF5F9",X"FFFAFE",X"FFF5F6",X"F9F7FA",X"F4F7FC",X"F4F9FC",X"F9F9F7",X"FEF6F3",X"FAEFEB",X"F6E8E5",X"FDF2E0",X"FDF1E1",X"FBF2E3",X"FAF2E5",X"FAF2E7",X"FAF2E7",X"F9F3E5",X"F9F3E5",X"FFF2EA",X"FFFCF3",X"FAFBF5",X"FFF7FC",X"F3F8FB",X"F0FBFD",X"FFFAFF",X"E7FAF8",X"F3F3F3",X"FAF9FE",X"F9EBFA",X"FCE2FB",X"F6EAFF",X"E6F0FC",X"EBEFFA",X"FAE8F8",X"FFE8F1",X"FFF7FB",X"FFF7F5",X"F8F7F3",X"F6F5F1",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FBFFFD",X"FFFEFB",X"F6EFF7",X"FAF7FF",X"FFFDFF",X"FCF8F7",X"F7FFFF",X"DBFFFF",X"F0F5FB",X"FFFDFF",X"F7FBFC",X"E6FCEF",X"E8FFF9",X"F8FFFF",X"EDF0F9",X"F6FFFC",X"EDFFFF",X"F4FFFF",X"FBFEFF",X"FBFBFB",X"FEFEFE",X"FBFBFD",X"FFFDFE",X"FFFBFC",X"FFFAFF",X"FFFCFF",X"F7F8FD",X"FFF0F5",X"FFECF3",X"FFF0F2",X"F8F6F9",X"FFF9FF",X"F9FBF6",X"FCFBF6",X"F5F5EB",X"FAFDF6",X"FBFFFF",X"F8FDFF",X"FEFFFF",X"FFFEF8",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFAFD",X"FBFFFA",X"F0FFF6",X"FFEDF1",X"F8E0F0",X"EFF3FF",X"FDF7FF",X"FFF2F9",X"FDEFFC",X"EFFCF5",X"FAEFFD",X"FCF3F8",X"F2FBFA",X"F1FBFD",X"E6F7ED",X"FFFDFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFD",X"FFFFF8",X"FFFDFF",X"FEFFFF",X"FEFFFB",X"FDFEFF",X"FEFFF2",X"FDFAFF",X"FFFCF8",X"F6FFF4",X"F7FEFF",X"FFF9FF",X"FFF8FF",X"F9FFF6",X"E7F1E9",X"FFFEFB",X"FFF4F7",X"FFF6F7",X"EFFFFE",X"FFFDFF",X"FFFCFA",X"F8FFF6",X"F6F9F0",X"F3F8F2",X"FCF1F9",X"FFFCFF",X"FFF7FA",X"FFF4FB",X"FFFAFF",X"F7FFFF",X"F9FFFF",X"FFFDFB",X"F5FFFB",X"F8FEFA",X"FFF5F4",X"F9EDDF",X"F7E6CC",X"ECE5BB",X"E0EAB6",X"FCDFB7",X"DCD1B1",X"DCDFB2",X"E9DBAA",X"F0D9A5",X"E5DFA5",X"D8D0A1",X"E7D6B8",X"BDC0A3",X"ABBBB0",X"C7ACB1",X"E2A8BE",X"E1A9C2",X"D4A6C0",X"DDA7C7",X"E8ABCD",X"E5A8CA",X"CAAEC4",X"B5AFB1",X"A5AEA9",X"9ED6CB",X"B6DAD6",X"A4D9C5",X"A9B2AD",X"C6AEBE",X"B5AFC9",X"D0A4C5",X"C7AFC5",X"BAB3C5",X"CAADC9",X"B8B0BF",X"9FAEA7",X"C2AFA8",X"D4ADB0",X"CAACB6",X"C1B1BC",X"B9AFB7",X"B7B1B3",X"A9ADAC",X"ACC4C8",X"A8CEDB",X"A2D2D4",X"BEC2C5",X"ADAAA3",X"A8BAAA",X"B0A6A4",X"D7A6A9",X"E4B9A8",X"E9C39F",X"E5B994",X"D9B792",X"ECC8A6",X"EEBBA0",X"DFAB96",X"E1C2B0",X"C0B1AA",X"B6AAAE",X"A8ABA0",X"ACA9A4",X"A99EA2",X"B5AAB2",X"A9A2AA",X"A8A6AB",X"A4A2A3",X"B8B4B3",X"C2ACA1",X"B1A8A3",X"C2B5AD",X"E9C5B5",X"EABDA8",X"E0C1AC",X"D6C1A2",X"DFC499",X"E9BC9D",X"EABEA1",X"E7BFA5",X"E1BFA6",X"DCBEA4",X"DABCA0",X"E9C4A7",X"EDC1A4",X"BDB7B7",X"BDB0B7",X"C1ADB8",X"B4A9B1",X"D8A9B9",X"CCB3B9",X"DDB9C5",X"DFA9C0",X"CAB4B7",X"FFF1FC"),
(X"FCFEFD",X"FFFBFD",X"F9FFFD",X"FFFBFF",X"E3FFFD",X"FFFDFF",X"F1FFFE",X"F2FFFB",X"F7FFFF",X"FAFDF6",X"FFFBF6",X"FFF3F9",X"FFF5FF",X"FFF6FF",X"FFF8FF",X"FBFFF9",X"FFF6FF",X"FFF9FF",X"FFF3FF",X"FFFAFF",X"FFFEF4",X"FFFEDB",X"FFFBE8",X"FFF9FF",X"F9FDFF",X"FFF9FF",X"FFF7FF",X"FFFCFF",X"FBFFFF",X"FFFBFF",X"FFFAFB",X"FFF7E9",X"FFFBF2",X"FFFDF1",X"FFF6F9",X"FFFAFF",X"FFFCED",X"F7FAEF",X"FFFDFF",X"FFFAFF",X"FFFCFF",X"FFF6FF",X"FFFAFF",X"FFFAFF",X"F9FDFF",X"FFFBFF",X"FFF5FF",X"FFFCE8",X"FFFFF3",X"FEF3ED",X"FFFFF4",X"F7FDF3",X"FFF7F9",X"FFFAF3",X"FFFFED",X"FEFEF6",X"FFFFF3",X"FFF6F6",X"FFFAF9",X"FFFBED",X"FBF9EA",X"FFFBFB",X"FFF0F4",X"F8FFF1",X"FFFEEA",X"FFFDED",X"FFFDF4",X"FFF8F8",X"FFF7FB",X"FFFCFF",X"FFFAFE",X"FFFAFE",X"FFFCFD",X"FFFEFF",X"FCFFFF",X"F8FDFF",X"FBFBF9",X"FFFAF7",X"FFFCF8",X"FFFBF8",X"FFFDEB",X"FFFDED",X"FFFEEF",X"FFFCEF",X"FFFCF1",X"FFFEF3",X"FFFFF1",X"FFFDEF",X"FFFAF2",X"FFFFF6",X"FBFCF6",X"FFF3F8",X"FBFFFF",X"F7FFFF",X"FFF2FB",X"F2FFFF",X"FCFCFC",X"FFFEFF",X"FFF4FF",X"FFF2FF",X"FFF9FF",X"F1FBFF",X"F8FCFF",X"FFF8FF",X"FFF6FF",X"FFF6FA",X"FFFAF8",X"FFFEFA",X"FFFFFB",X"FFFDFE",X"F9F7FC",X"FDFCFF",X"FBFFFD",X"F6F2EF",X"FFFCFF",X"FCF9FF",X"FFFCFF",X"FCF8F7",X"F7FFFF",X"E1FFFF",X"F8FDFF",X"FFFCFF",X"F8FCFD",X"F1FFFA",X"ECFFFD",X"F4FCFF",X"FCFFFF",X"F5FFFB",X"EEFFFF",X"EEFAFF",X"FCFFFF",X"FCFCFC",X"FFFFFF",X"FEFEFF",X"FFFDFE",X"FFFEFF",X"FFF9FF",X"FFFDFF",X"FBFCFF",X"FFF9FE",X"FFF1F8",X"FFF3F5",X"FFFEFF",X"FFFBFF",X"FCFEF9",X"FBFAF5",X"FFFFF6",X"FBFEF7",X"FCFFFF",X"FBFFFF",X"FEFFFF",X"FFFDF7",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFAFD",X"F9FFF8",X"EEFFF4",X"FFF7FB",X"FFF6FF",X"F5F9FF",X"FFFBFF",X"FFF7FE",X"FFF7FF",X"F7FFFD",X"FFFAFF",X"FFF8FD",X"F9FFFF",X"F8FFFF",X"F3FFFA",X"FAF8FF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFD",X"FFFFF8",X"FFFDFF",X"FEFFFF",X"FEFFFB",X"FDFEFF",X"FEFFF2",X"FDFAFF",X"FFFEFA",X"F5FFF3",X"F8FFFF",X"FFF8FF",X"FFFAFF",X"F4FFF1",X"F9FFFB",X"FDF8F5",X"FFF7FA",X"FFF8F9",X"F2FFFF",X"FFFAFC",X"FFF7F5",X"F8FFF6",X"FDFFF7",X"FBFFFA",X"FFFAFF",X"FDF8FC",X"FFFCFF",X"FFF9FF",X"FFFDFF",X"F7FFFF",X"EFF8F5",X"FFFDFB",X"F7FFFD",X"F6FCF8",X"FFFBFA",X"FFFDEF",X"FFFAE0",X"FFFFD8",X"F9FFCF",X"FFF9D1",X"FFFFDF",X"FFFFD6",X"FFFDCC",X"FFF9C5",X"FFFFCA",X"FFFFD2",X"FFFDDF",X"FFFFE5",X"F5FFFA",X"FFF5FA",X"FFE9FF",X"FFEAFF",X"FFEBFF",X"FFE7FF",X"FFE5FF",X"FFE4FF",X"FFF3FF",X"FEF8FA",X"F9FFFD",X"D4FFFF",X"E6FFFF",X"D6FFF7",X"F9FFFD",X"FFF0FF",X"FFFAFF",X"FFEEFF",X"FFF1FF",X"FEF7FF",X"FFF3FF",X"FFFAFF",X"F5FFFD",X"FFFAF3",X"FFEFF2",X"FFF3FD",X"FFF9FF",X"FFF8FF",X"FFFDFF",X"FCFFFF",X"EBFFFF",X"E1FFFF",X"D8FFFF",X"F8FCFF",X"FFFFF8",X"EEFFF0",X"FFFCFA",X"FFF0F3",X"FFF4E3",X"FFF3CF",X"FFF4CF",X"FFF7D2",X"FFF0CE",X"FFF0D5",X"FFF2DD",X"FFF6E4",X"FFF6EF",X"FFFBFF",X"FCFFF4",X"FFFFFA",X"FFFBFF",X"FFF5FD",X"FFFCFF",X"FFFDFF",X"FFFEFF",X"FFFBFA",X"FFF9EE",X"FFFDF8",X"FFF7EF",X"FFF6E6",X"FFF2DD",X"FFF4DF",X"FFF8D9",X"FFFCD1",X"FFF3D4",X"FFF2D5",X"FFF2D8",X"FFF8DF",X"FFF6DC",X"FFF9DD",X"FFF4D7",X"FFF5D8",X"FFFCFC",X"FFF7FE",X"FFF8FF",X"FFFBFF",X"FFEAFA",X"FFF6FC",X"FFF2FE",X"FFE7FE",X"FFF8FB",X"FFF5FF"),
(X"FFFDFF",X"FEFFFF",X"FCFFFF",X"FFFFFD",X"FFFDFD",X"FFFBFF",X"FFFEFF",X"FEFFFF",X"FBFDFF",X"FDFFFE",X"FEFFFA",X"FFFBFF",X"FFFBFF",X"FFFFFD",X"FEFFFA",X"FCFFFF",X"FFFEFB",X"FFFEFD",X"FFFEFF",X"FFFDFF",X"FFFEFF",X"FFFEFF",X"FFFFFD",X"FFFFFB",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFB",X"FCFFFB",X"FEFFFB",X"FEFFFD",X"FFFFFF",X"FFFEFF",X"FBFFFB",X"FCFFFA",X"FEFFF8",X"FFFFF8",X"FFFFFA",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FEFFFD",X"FEFFFD",X"FFFFFB",X"FFFFFB",X"FFFFFD",X"FFFEFF",X"FFFEFF",X"FFFDFF",X"FEFFFF",X"FFFEFF",X"FFFDFD",X"FFFDFB",X"FFFEFD",X"FFFFFD",X"FFFFFA",X"FFFEF8",X"FFFEFF",X"FFFEFF",X"FFFFFD",X"FFFFFD",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFD",X"FCFFFB",X"FCFFFB",X"FFFFFF",X"FFFDFF",X"FFFDFF",X"FEFFFD",X"F9FFF8",X"FFFEFF",X"FEFFFF",X"FCFFFB",X"FEFFFD",X"FFFEFF",X"FFFDFF",X"FFFFFD",X"FFFFFA",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FCFFFB",X"FFFFFD",X"FFFDFF",X"FFFEFF",X"FCFFFF",X"F9FFFF",X"FEFFFD",X"FFFEFB",X"F9FFFD",X"FEFFFD",X"FFFFFD",X"FFFFFD",X"FEFFFD",X"FCFFFD",X"FEFFFD",X"FFFEFD",X"FFFCFF",X"FFFFFF",X"FBFFFF",X"FBFFFF",X"FEFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FEFFFF",X"F9FFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFFFD",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFD",X"FFFFFD",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFB",X"FFFEFB",X"FFFFFF",X"FBFFFF",X"FCFFFF",X"FFFFFF",X"FFFDFF",X"FFFEFF",X"FFFFFF",X"FCFFFF",X"FCFFFF",X"FEFFFF",X"FFFFFD",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FEFFFF",X"FBFFFD",X"F9FFFD",X"F7FFFF",X"FFFBFF",X"FFF9FF",X"FEFFFF",X"F9FFFD",X"FFFFFD",X"FFFEFB",X"FCFFFB",X"FFFEF8",X"FEFFFF",X"F9FFFF",X"F9FFFF",X"FFFFFB",X"FFFFF8",X"FFFFFB",X"FCFFFF",X"FFFDFB",X"FFFEFB",X"FFFFFF",X"FFFDFF",X"FFFAFF",X"FFFAFF",X"FFFFFF",X"F8FFFA",X"FFFDFF",X"FFFFFF",X"FEFFFD",X"FFFFFB",X"FFFFFA",X"FFFEFB",X"FFFEFD",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFD",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFF8",X"FFFFF3",X"FFFFFD",X"FFFDFF",X"FFFEFF",X"FEFFF8",X"FEFFF3",X"FEFFFB",X"FFFFFF",X"FFFFFB",X"FCFFFD",X"FEFFFF",X"FFFFFF",X"FFFDFF",X"FFFDFF",X"FFFEFF",X"FFFFFF",X"FEFFFD",X"FFFDFB",X"FFFFFD",X"FCFFFF",X"FBFFFF",X"FCFFFF",X"FEFFFF",X"FCFFFF",X"FBFFFF",X"FEFFFF",X"FFFFFF",X"FFFDFF",X"FFFCFF",X"FFFCFF",X"FFFDFF",X"FFFEFF",X"FCFFFF",X"FDFEFF",X"FBFFFF",X"FAFFFE",X"F8FFFE",X"F8FFFE",X"FAFFFE",X"FBFFFF",X"FDFEFF",X"FCFEF9",X"FCFEFD",X"FDFDFF",X"FDFDFD",X"FDFEF9",X"FCFFF8",X"FAFFF9",X"FAFEFD",X"FDFFFA",X"FDFFFA",X"FDFFFA",X"FDFFFA",X"FEFFFA",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"F7FFFE",X"FBFFFE",X"FFFDFE",X"FFFDFE",X"FDFFFE",X"FBFFFE",X"FDFFFE",X"FFFDFE",X"FEFEFE",X"FBFFFE",X"FBFFFE",X"FDFFFE",X"FFFDFE",X"FFFBFE",X"FFFCFE",X"FFFDFE",X"FFFDFC",X"FFFEFC",X"FEFEFC",X"FDFFFE",X"FDFFFE",X"FBFFFF",X"FBFFFF",X"FBFFFF",X"FDFFFE",X"FDFFFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFFFF",X"FFFFFF",X"FFFDFF",X"FFFBFF",X"FFFCFF",X"FFFDFF",X"FFFFFF",X"FEFFFD",X"F6FFFE",X"FDFFFE",X"FFFBFE",X"FFFBFF",X"FEFEFF",X"F8FFFF",X"F8FFFF",X"FAFFFF",X"FFFAFF",X"FFFDFF",X"FAFFFF",X"FBFFFF",X"FFFDFF",X"FFFBFF",X"FFFCFF",X"FEFDFF",X"FBFFFC",X"FDFFFC",X"FFFDFE",X"FEFEFE",X"FAFFFE",X"F8FFFE",X"F8FFFE",X"FAFFFE",X"FDFFFE",X"FDFFFE"),
(X"FFFDFF",X"FEFFFF",X"FCFFFF",X"FFFFFD",X"FFFDFD",X"FFFBFF",X"FFFEFF",X"FEFFFF",X"FBFDFF",X"FDFFFE",X"FEFFFA",X"FFFBFF",X"FFFCFF",X"FFFFFD",X"FEFFFA",X"FCFFFF",X"FFFEFB",X"FFFEFD",X"FFFEFF",X"FFFDFF",X"FFFEFF",X"FFFEFF",X"FFFFFD",X"FFFFFB",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFB",X"FCFFFB",X"FEFFFB",X"FEFFFD",X"FFFFFF",X"FFFEFF",X"FBFFFB",X"FCFFFA",X"FEFFF8",X"FFFFF8",X"FFFFFA",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FEFFFD",X"FEFFFD",X"FFFFFB",X"FFFFFB",X"FFFFFD",X"FFFEFF",X"FFFEFF",X"FFFDFF",X"FEFFFF",X"FFFEFF",X"FFFDFD",X"FFFDFB",X"FFFEFD",X"FFFFFD",X"FFFFFA",X"FFFEF8",X"FFFEFF",X"FFFEFF",X"FFFFFD",X"FFFFFD",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFD",X"FCFFFB",X"FCFFFB",X"FFFFFF",X"FFFDFF",X"FFFDFF",X"FEFFFD",X"F9FFF8",X"FFFEFF",X"FEFFFF",X"FCFFFB",X"FEFFFD",X"FFFEFF",X"FFFDFF",X"FFFFFD",X"FFFFFA",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FCFFFB",X"FFFFFD",X"FFFDFF",X"FFFEFF",X"FCFFFF",X"F9FFFF",X"FEFFFD",X"FFFEFB",X"F9FFFD",X"FEFFFD",X"FFFFFD",X"FFFFFD",X"FEFFFD",X"FCFFFD",X"FEFFFD",X"FFFEFD",X"FFFCFF",X"FFFFFF",X"FBFFFF",X"FBFFFF",X"FEFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FEFFFF",X"F9FFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFFFD",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFD",X"FFFFFD",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFB",X"FFFEFB",X"FFFFFF",X"FBFFFF",X"FCFFFF",X"FFFFFF",X"FFFDFF",X"FFFEFF",X"FFFFFF",X"FCFFFF",X"FCFFFF",X"FEFFFF",X"FFFFFD",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FEFFFF",X"FBFFFD",X"F9FFFD",X"F7FFFF",X"FFFBFF",X"FFF9FF",X"FEFFFF",X"F9FFFD",X"FFFFFD",X"FFFEFB",X"FCFFFB",X"FFFEF8",X"FEFFFF",X"F9FFFF",X"F9FFFF",X"FFFFFB",X"FFFFF8",X"FFFFFB",X"FCFFFF",X"FFFDFB",X"FFFEFB",X"FFFFFF",X"FFFDFF",X"FFFAFF",X"FFFAFF",X"FFFFFF",X"F8FFFA",X"FFFDFF",X"FFFFFF",X"FEFFFD",X"FFFFFB",X"FFFFFA",X"FFFEFB",X"FFFEFD",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFD",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFF8",X"FFFFF3",X"FFFFFD",X"FFFDFF",X"FFFEFF",X"FEFFF8",X"FEFFF3",X"FEFFFB",X"FFFFFF",X"FFFFFB",X"FCFFFD",X"FEFFFF",X"FFFFFF",X"FFFDFF",X"FFFDFF",X"FFFEFF",X"FFFFFF",X"FEFFFD",X"FFFDFB",X"FFFFFD",X"FCFFFF",X"FBFFFF",X"FCFFFF",X"FEFFFF",X"FCFFFF",X"FBFFFF",X"FEFFFF",X"FFFFFF",X"FFFDFF",X"FFFCFF",X"FFFCFF",X"FFFDFF",X"FFFEFF",X"FCFFFF",X"FDFEFF",X"FBFFFF",X"FAFFFE",X"F8FFFE",X"F8FFFE",X"FAFFFE",X"FBFFFF",X"FDFEFF",X"FDFFFA",X"FDFFFE",X"FEFEFF",X"FEFEFE",X"FEFFFA",X"FDFFF9",X"FBFFFA",X"FBFFFE",X"FDFFFA",X"FDFFFA",X"FDFFFA",X"FDFFFA",X"FEFFFA",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"F7FFFE",X"FBFFFE",X"FFFDFE",X"FFFDFE",X"FDFFFE",X"FBFFFE",X"FDFFFE",X"FFFDFE",X"FEFEFE",X"FBFFFE",X"FBFFFE",X"FDFFFE",X"FFFDFE",X"FFFBFE",X"FFFCFE",X"FFFDFE",X"FFFDFC",X"FFFEFC",X"FEFEFC",X"FDFFFE",X"FDFFFE",X"FBFFFF",X"FBFFFF",X"FBFFFF",X"FDFFFE",X"FDFFFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FEFFFF",X"FFFFFF",X"FFFDFF",X"FFFBFF",X"FFFCFF",X"FFFDFF",X"FFFFFF",X"FEFFFD",X"F6FFFE",X"FDFFFE",X"FFFBFE",X"FFFBFF",X"FEFEFF",X"F8FFFF",X"F8FFFF",X"FAFFFF",X"FFFAFF",X"FFFDFF",X"FAFFFF",X"FBFFFF",X"FFFDFF",X"FFFBFF",X"FFFCFF",X"FEFDFF",X"FBFFFC",X"FDFFFC",X"FFFDFE",X"FEFEFE",X"FAFFFE",X"F8FFFE",X"F8FFFE",X"FAFFFE",X"FDFFFE",X"FDFFFE"),
(X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFD",X"FFFFFD",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FFFFFF",X"FFFFFD",X"FFFFFD",X"FFFEFF",X"FFFFFF",X"FFFFFB",X"FFFFFB",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FCFFFF",X"FCFFFF",X"FBFFFF",X"FBFFFF",X"FCFFFF",X"FCFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFAFF",X"FFFCFF",X"FFFEFF",X"FCFFFF",X"FBFFFF",X"FCFFFF",X"FFFFFF",X"FFFEFF",X"FFFDFF",X"FFFEFF",X"FFFEFF",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FEFFFD",X"FFFEFA",X"FFFEFF",X"FCFFFF",X"FCFFFF",X"FEFFFF",X"FEFFFF",X"FBFFFF",X"F8FFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFFFF",X"FEFFFD",X"FFFFFF",X"FFFEFF",X"FFFDFF",X"FFFFFF",X"FCFFFD",X"FFFDFF",X"FFFEFF",X"FFFFFD",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FCFFFD",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"F8FFFF",X"FCFFFF",X"FFFFFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FBFFFF",X"FBFFFF",X"FFFCFF",X"FFFEFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FEFFFF",X"F9FFFF",X"F7FFFF",X"FFFEFF",X"FFFFFF",X"FCFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFD",X"FFFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFB",X"FFFEFB",X"FFFFFD",X"FEFFFF",X"FCFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFD",X"FEFFFF",X"FFFCFF",X"FFFDFF",X"F5FFFF",X"F4FFFF",X"FEFFFF",X"FFFEFF",X"FCFFFF",X"FFFEFD",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FCFFFD",X"F8FFFB",X"F7FFFB",X"F8FFFD",X"FCFFFD",X"FEFFFB",X"FFFFF8",X"FFFDFF",X"FFFFFF",X"FCFFFF",X"FCFFFF",X"FFFFFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFA",X"FFFFFA",X"FFFFFD",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFFEF",X"FFFFFA",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFDFF",X"FFFCFF",X"FFFDFF",X"FFFEFD",X"FFFFFF",X"FCFFFF",X"FBFFFF",X"FBFFFF",X"FEFFFF",X"FFFEFF",X"FFFEFD",X"FFFFFD",X"FEFFFF",X"FCFFFF",X"FEFFFF",X"FFFEFF",X"FFFDFF",X"FFFEFF",X"FFFFFD",X"FFFCFF",X"FFFFFF",X"F9FFFF",X"FBFFFF",X"FFFEFF",X"FFFDFF",X"FFFEFF",X"FBFFFF",X"FFFDFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFDFF",X"FEFFFD",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFB",X"FEFFFB",X"FEFFFF",X"FEFFFF",X"FFFCFF",X"FFFDFF",X"FFFEFF",X"FFFFFB",X"FFFFFF",X"FFFDFF",X"FEFFFF",X"FEFFF6",X"FCFFFF",X"FFFEFF",X"FFFDFF",X"FFFCFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFFFF",X"FCFFFF",X"FFFFFD",X"FFFFFD",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFDFF",X"FFFDFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFFFF",X"FCFFFA",X"FCFFF8",X"FCFFF8",X"FCFFFA",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FCFFFF",X"FEFFFF",X"FFFFFF",X"FFFDFF",X"F4FFFF",X"F7FFFF",X"F9FFFF",X"FEFFFF",X"FFFEFF",X"FFFEFF",X"FEFFFF",X"FBFFFF",X"FCFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FFFEFF",X"FFFDFF",X"FFFFFF",X"FFFFFF"),
(X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFD",X"FFFFFD",X"FFFDFE",X"FEFEFE",X"FDFEFF",X"FFFFFF",X"FFFFFD",X"FFFFFD",X"FFFEFF",X"FFFFFF",X"FFFFFB",X"FFFFFB",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FCFFFF",X"FCFFFF",X"FBFFFF",X"FBFFFF",X"FCFFFF",X"FCFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFAFF",X"FFFCFF",X"FFFEFF",X"FCFFFF",X"FBFFFF",X"FCFFFF",X"FFFFFF",X"FFFEFF",X"FFFDFF",X"FFFEFF",X"FFFEFF",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FEFFFD",X"FFFEFA",X"FFFEFF",X"FCFFFF",X"FCFFFF",X"FEFFFF",X"FEFFFF",X"FBFFFF",X"F8FFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFFFF",X"FEFFFD",X"FFFFFF",X"FFFEFF",X"FFFDFF",X"FFFFFF",X"FCFFFD",X"FFFDFF",X"FFFEFF",X"FFFFFD",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FCFFFD",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"F8FFFF",X"FCFFFF",X"FFFFFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FBFFFF",X"FBFFFF",X"FFFCFF",X"FFFEFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FEFFFF",X"F9FFFF",X"F7FFFF",X"FFFEFF",X"FFFFFF",X"FCFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFD",X"FFFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFB",X"FFFEFB",X"FFFFFD",X"FEFFFF",X"FCFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFD",X"FEFFFF",X"FFFCFF",X"FFFDFF",X"F5FFFF",X"F4FFFF",X"FEFFFF",X"FFFEFF",X"FCFFFF",X"FFFEFD",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FCFFFD",X"F8FFFB",X"F7FFFB",X"F8FFFD",X"FCFFFD",X"FEFFFB",X"FFFFF8",X"FFFDFF",X"FFFFFF",X"FCFFFF",X"FCFFFF",X"FFFFFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFA",X"FFFFFA",X"FFFFFD",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFFEF",X"FFFFFA",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFDFF",X"FFFCFF",X"FFFDFF",X"FFFEFD",X"FFFFFF",X"FCFFFF",X"FBFFFF",X"FBFFFF",X"FEFFFF",X"FFFEFF",X"FFFEFD",X"FFFFFD",X"FEFFFF",X"FCFFFF",X"FEFFFF",X"FFFEFF",X"FFFDFF",X"FFFEFF",X"FFFFFD",X"FFFCFF",X"FFFFFF",X"F9FFFF",X"FBFFFF",X"FFFEFF",X"FFFDFF",X"FFFEFF",X"FBFFFF",X"FFFDFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFDFF",X"FEFFFD",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFB",X"FEFFFB",X"FEFFFF",X"FEFFFF",X"FFFCFF",X"FFFDFF",X"FFFEFF",X"FFFFFB",X"FFFFFF",X"FFFDFF",X"FEFFFF",X"FEFFF6",X"FCFFFF",X"FFFEFF",X"FFFDFF",X"FFFCFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFFFF",X"FCFFFF",X"FFFFFD",X"FFFFFD",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFDFF",X"FFFDFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFFFF",X"FCFFFA",X"FCFFF8",X"FCFFF8",X"FCFFFA",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FCFFFF",X"FEFFFF",X"FFFFFF",X"FFFDFF",X"F4FFFF",X"F7FFFF",X"F9FFFF",X"FEFFFF",X"FFFEFF",X"FFFEFF",X"FEFFFF",X"FBFFFF",X"FCFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FFFEFF",X"FFFDFF",X"FFFFFF",X"FFFFFF"),
(X"FCFFFF",X"FFFFFF",X"FFFEFD",X"FFFFFD",X"FCFFFD",X"FAFFFE",X"FBFFFF",X"FEFCFF",X"FFFDF9",X"FFFCFF",X"FFFEFF",X"FEFFFD",X"FEFFF8",X"FFFFFA",X"FFFEFF",X"FFFDFF",X"FFFDFF",X"FFFEFF",X"FEFFFF",X"FCFFFF",X"FCFFFF",X"FCFFFF",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFD",X"FEFFFD",X"FEFFFD",X"FFFFFF",X"FFFEFF",X"FFFDFF",X"FFFCFF",X"FFFCFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FCFFFF",X"FEFFFF",X"FFFEFF",X"FFFDFF",X"FFFDFF",X"FFFDFF",X"FFFEFD",X"FFFEFB",X"FFFDFF",X"FFFDFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FEFFFB",X"FEFFFA",X"FCFFF8",X"FFFFF6",X"FFFFFD",X"F9FFFF",X"FBFFFF",X"FFFFFF",X"FFFFFB",X"FFFFFD",X"FBFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFD",X"FFFFFD",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFDFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FFFEFF",X"FEFFFF",X"FCFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFBFF",X"FFFEFF",X"F9FFFF",X"F8FFFF",X"FCFFFF",X"FFFEFF",X"FFFDFF",X"FFFEFF",X"FFFDFF",X"FFFDFF",X"FFFDFF",X"FFFDFF",X"FFFBFF",X"FFFAFF",X"FFFBFF",X"FFFBFF",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFD",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FFFFFD",X"FFFFFB",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FFFEFD",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FFFFFF",X"FFFFFD",X"FFFFFD",X"FFFFFB",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFDFF",X"FFFDFF",X"FFFEFF",X"FFFEFF",X"FEFFFF",X"F8FFFF",X"FBFFFF",X"FFFDFF",X"FFFCFF",X"F9FFFF",X"FFFDFF",X"FFFBFF",X"FFFBFB",X"FFFBFD",X"FFFCFF",X"FFFDFF",X"FFFCFF",X"FFFBFD",X"FFFDFF",X"FFFDFF",X"FFFCFD",X"FFFEF8",X"FFFFF6",X"FFFFF8",X"FFFCFB",X"FFF9FD",X"FFFEFD",X"FFFFFF",X"FCFFFF",X"FBFFFF",X"FBFFFF",X"FCFFFF",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFD",X"FFFFFA",X"FFFFFB",X"FFFEFF",X"FEFDFF",X"FEFCFF",X"FEFCFF",X"FFFDFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFF8",X"FFFFF6",X"FFFFF8",X"FFFDFF",X"FFFCFF",X"FFFCFD",X"FFFCFB",X"FFFCFB",X"FFFCFD",X"FFFDFF",X"FFFEFF",X"FCFFFF",X"FCFFFF",X"FFFFFF",X"FFFEFF",X"FFFDFF",X"FFFDFF",X"FFFDFD",X"FFFEFB",X"FFFBFF",X"FEFFFF",X"F5FFFF",X"F7FFFF",X"FEFFFF",X"FFFDFF",X"FFFEFF",X"FBFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFDFF",X"FFFDFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFCFF",X"FFFCFF",X"FFFDFF",X"FFFFF6",X"FFFFFF",X"FFFCFF",X"FEFEFF",X"FEFFF1",X"FFFDFF",X"FFFEFF",X"FFFEFF",X"FEFFFF",X"FCFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FCFFFF",X"FCFFFF",X"FBFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFDFF",X"FFFDFF",X"FFFDFF",X"FFFCFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFDFF",X"FFFFFF",X"FBFFFB",X"F8FFFA",X"F8FFFA",X"FBFFFD",X"FFFFFF",X"FFFDFF",X"FFFBFF",X"FFFEFF",X"F9FFFF",X"F8FFFF",X"FCFFFF",X"FFFEFF",X"FFFDFF",X"FFFDFF",X"F7FFFD",X"FCFFFD",X"FFFFFD",X"FFFFFD",X"FCFFFD",X"FBFFFB",X"FCFFFB",X"FFFFFB",X"FFFEFF",X"FFFDFF",X"FFFBFF",X"FFFBFF",X"FFFCFF",X"FFFCFF",X"FFFBFF",X"FFF9FF",X"FFFFFF",X"FFFEFF"),
(X"FCFFFF",X"FFFFFF",X"FFFEFD",X"FFFFFD",X"FCFFFD",X"FAFFFE",X"FAFEFF",X"FDFBFF",X"FFFCF8",X"FFFBFF",X"FEFDFF",X"FEFFFD",X"FEFFF8",X"FFFFFA",X"FFFEFF",X"FFFDFF",X"FFFDFF",X"FFFEFF",X"FEFFFF",X"FCFFFF",X"FCFFFF",X"FCFFFF",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFD",X"FEFFFD",X"FEFFFD",X"FFFFFF",X"FFFEFF",X"FFFDFF",X"FFFCFF",X"FFFCFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FCFFFF",X"FEFFFF",X"FFFEFF",X"FFFDFF",X"FFFDFF",X"FFFDFF",X"FFFEFD",X"FFFEFB",X"FFFDFF",X"FFFDFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FEFFFB",X"FEFFFA",X"FCFFF8",X"FFFFF6",X"FFFFFD",X"F9FFFF",X"FBFFFF",X"FFFFFF",X"FFFFFB",X"FFFFFD",X"FBFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFD",X"FFFFFD",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFDFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FFFEFF",X"FEFFFF",X"FCFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFBFF",X"FFFEFF",X"F9FFFF",X"F8FFFF",X"FCFFFF",X"FFFEFF",X"FFFDFF",X"FFFEFF",X"FFFDFF",X"FFFDFF",X"FFFDFF",X"FFFDFF",X"FFFBFF",X"FFFAFF",X"FFFBFF",X"FFFBFF",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFD",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FFFFFD",X"FFFFFB",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FFFEFD",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FFFFFF",X"FFFFFD",X"FFFFFD",X"FFFFFB",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFDFF",X"FFFDFF",X"FFFEFF",X"FFFEFF",X"FEFFFF",X"F8FFFF",X"FBFFFF",X"FFFDFF",X"FFFCFF",X"F9FFFF",X"FFFDFF",X"FFFBFF",X"FFFBFB",X"FFFBFD",X"FFFCFF",X"FFFDFF",X"FFFCFF",X"FFFBFD",X"FFFDFF",X"FFFDFF",X"FFFCFD",X"FFFEF8",X"FFFFF6",X"FFFFF8",X"FFFCFB",X"FFF9FD",X"FFFEFD",X"FFFFFF",X"FCFFFF",X"FBFFFF",X"FBFFFF",X"FCFFFF",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFD",X"FFFFFA",X"FFFFFB",X"FFFEFF",X"FEFDFF",X"FEFCFF",X"FEFCFF",X"FFFDFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFF8",X"FFFFF6",X"FFFFF8",X"FFFDFF",X"FFFCFF",X"FFFCFD",X"FFFCFB",X"FFFCFB",X"FFFCFD",X"FFFDFF",X"FFFEFF",X"FCFFFF",X"FCFFFF",X"FFFFFF",X"FFFEFF",X"FFFDFF",X"FFFDFF",X"FFFDFD",X"FFFEFB",X"FFFBFF",X"FEFFFF",X"F5FFFF",X"F7FFFF",X"FEFFFF",X"FFFDFF",X"FFFEFF",X"FBFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFDFF",X"FFFDFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FEFEFF",X"FEFEFE",X"FEFEFC",X"FEFEFC",X"FEFEFC",X"FEFEFE",X"FEFDFF",X"FEFDFF",X"FFFCFF",X"FFFCFF",X"FFFDFF",X"FFFFF6",X"FFFFFF",X"FFFCFF",X"FEFEFF",X"FEFFF1",X"FFFDFF",X"FFFEFF",X"FFFEFF",X"FEFFFF",X"FCFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FCFFFF",X"FCFFFF",X"FBFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFDFF",X"FFFDFF",X"FFFDFF",X"FFFCFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFDFF",X"FFFFFF",X"FBFFFB",X"F8FFFA",X"F8FFFA",X"FBFFFD",X"FFFFFF",X"FFFDFF",X"FFFBFF",X"FFFEFF",X"F9FFFF",X"F8FFFF",X"FCFFFF",X"FFFEFF",X"FFFDFF",X"FFFDFF",X"F7FFFD",X"FCFFFD",X"FFFFFD",X"FFFFFD",X"FCFFFD",X"FBFFFB",X"FCFFFB",X"FFFFFB",X"FFFEFF",X"FFFDFF",X"FFFBFF",X"FFFBFF",X"FFFCFF",X"FFFCFF",X"FFFBFF",X"FFF9FF",X"FFFFFF",X"FFFEFF"),
(X"FBFFFE",X"FFFEFF",X"FFFCFD",X"FFFEFD",X"FCFFFF",X"FAFFFF",X"FDFCFF",X"FFF7FF",X"FFF5FF",X"FFF7FF",X"FEFAFF",X"FDFFFE",X"FCFFF8",X"FEFFFB",X"FFFDFF",X"FFFCFF",X"FFFAFF",X"FFFBFF",X"FFFDFD",X"FFFEFB",X"FFFFFB",X"FFFEFD",X"FFFDFF",X"FFFCFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFD",X"FEFFFD",X"FEFFFD",X"FEFFFD",X"FCFFFD",X"FEFFFF",X"FFFEFF",X"FFFDFF",X"FFFDFF",X"FFFEFF",X"FEFFFB",X"FBFFFA",X"FEFFFB",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FCFFFF",X"FCFFFF",X"FCFFFD",X"FCFFFB",X"FEFFFD",X"FEFFFF",X"FEFFFF",X"FCFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFD",X"FFFFFB",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFD",X"FFFDF8",X"FFFCF3",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFD",X"FFFFFD",X"FFFFFB",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFFFD",X"FCFFFB",X"FCFFFD",X"FFFFFF",X"FFFDFF",X"FCFFFB",X"FEFFFD",X"FFFFFF",X"FFFFFF",X"FEFFFD",X"FEFFFD",X"FEFFFF",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFF9FF",X"FFFEFF",X"F9FFFD",X"F9FFFB",X"FFFFFB",X"FFFCFD",X"FFFDFF",X"FFFEFF",X"F8FFFF",X"FCFFFF",X"FFFFFF",X"FEFFFF",X"F9FFFF",X"F9FFFF",X"FEFFFF",X"FFFDFF",X"FBFFFF",X"FEFFFF",X"FFFEFF",X"FFFDFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FCFFFF",X"FEFFFF",X"FEFFFF",X"FCFFFF",X"FBFFFF",X"FCFFFF",X"FFFFFF",X"FFFEFF",X"FFFFFD",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FFFFFB",X"FFFFFA",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFFFD",X"FFFFFD",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FCFFFF",X"FCFFFF",X"FFFFFF",X"FFFEFD",X"FFFEFF",X"FEFFFF",X"FCFFFF",X"FCFFFF",X"FEFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFCFF",X"FFFDFF",X"FFFFFF",X"FEFFFF",X"FCFFFD",X"FCFFFD",X"FEFFFD",X"FEFFFD",X"FEFFFB",X"FCFFFB",X"FCFFFD",X"FFFFFD",X"FFFBFF",X"FFF9FF",X"FFFDFF",X"F9FFFF",X"F4FFFF",X"FBFFFF",X"FFFFF8",X"FFFFFA",X"F8FFFF",X"F5FFFF",X"F8FFFF",X"FCFFFA",X"F1FFFF",X"F9FFFF",X"FFFDFF",X"FFFDFF",X"FCFFFF",X"F8FFFF",X"F9FFFF",X"FEFFFF",X"FFFFFB",X"FFFFFD",X"FFFEFF",X"FEFFFF",X"FCFFFF",X"FCFFFF",X"FFFFFF",X"FFFEFD",X"FEFFFF",X"FFFFFF",X"FFFFFB",X"FFFFFA",X"FFFFFB",X"FEFFFA",X"FEFFF4",X"FCFFF1",X"FEFEFF",X"FEFFFA",X"FEFFF3",X"FFFFF6",X"FFFFF8",X"FFFFF8",X"FFFFFD",X"FEFFFF",X"FFFDFF",X"FFFFFF",X"F9FFFB",X"F5FFFA",X"F5FFFA",X"F8FFFB",X"FCFFFF",X"FFFEFF",X"FBFFFF",X"FEFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFD",X"FFFFFD",X"FFFFFB",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFD",X"FEFFFD",X"F9FFFD",X"FBFFFD",X"FCFFFF",X"FEFFFF",X"FEFFFF",X"FCFFFF",X"FBFFFD",X"F9FFFD",X"FFFEFF",X"FFFFFF",X"FFFFFB",X"FFFFFB",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFF1",X"FFFFFF",X"FFFFFF",X"FFFFF4",X"FFFFF6",X"FFFDFF",X"FFFDFF",X"FFFFF6",X"FFFBFF",X"FFFEFF",X"FBFFFF",X"F8FFFF",X"F9FFFF",X"FCFFFF",X"FEFFFF",X"FFFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FCFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFD",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFDFF",X"FFFEFF",X"FFFEFF",X"FFFAFF",X"FFFEFF",X"F9FFFF",X"F9FFFF",X"FFFFFF",X"FFFEFF",X"FFFFFF",X"FBFFFF",X"FFFBFF",X"FFFAFF",X"FFFAFF",X"FFFEFD",X"F9FFFD",X"F8FFFD",X"FEFFFB",X"FFFDFB",X"F8FFFF",X"F9FFFF",X"FBFFFF",X"F9FFFF",X"F7FFFF",X"F7FFFF",X"F9FFFF",X"FCFFFF",X"FEFFFF",X"FEFFFF"),
(X"FBFFFE",X"FFFEFF",X"FFFCFD",X"FFFEFD",X"FCFFFF",X"FAFFFF",X"FCFBFF",X"FFF7FF",X"FFF4FE",X"FFF6FF",X"FEFAFF",X"FDFFFE",X"FCFFF8",X"FEFFFB",X"FFFDFF",X"FFFCFF",X"FFFAFF",X"FFFBFF",X"FFFDFD",X"FFFEFB",X"FFFFFB",X"FFFEFD",X"FFFDFF",X"FFFCFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFD",X"FEFFFD",X"FEFFFD",X"FEFFFD",X"FCFFFD",X"FEFFFF",X"FFFEFF",X"FFFDFF",X"FFFDFF",X"FFFEFF",X"FEFFFB",X"FBFFFA",X"FEFFFB",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FCFFFF",X"FCFFFF",X"FCFFFD",X"FCFFFB",X"FEFFFD",X"FEFFFF",X"FEFFFF",X"FCFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFD",X"FFFFFB",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFD",X"FFFDF8",X"FFFCF3",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFD",X"FFFFFD",X"FFFFFB",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFFFD",X"FCFFFB",X"FCFFFD",X"FFFFFF",X"FFFDFF",X"FCFFFB",X"FEFFFD",X"FFFFFF",X"FFFFFF",X"FEFFFD",X"FEFFFD",X"FEFFFF",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFF9FF",X"FFFEFF",X"F9FFFD",X"F9FFFB",X"FFFFFB",X"FFFCFD",X"FFFDFF",X"FFFEFF",X"F8FFFF",X"FCFFFF",X"FFFFFF",X"FEFFFF",X"F9FFFF",X"F9FFFF",X"FEFFFF",X"FFFDFF",X"FBFFFF",X"FEFFFF",X"FFFEFF",X"FFFDFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FCFFFF",X"FEFFFF",X"FEFFFF",X"FCFFFF",X"FBFFFF",X"FCFFFF",X"FFFFFF",X"FFFEFF",X"FFFFFD",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FFFFFB",X"FFFFFA",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFFFD",X"FFFFFD",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FCFFFF",X"FCFFFF",X"FFFFFF",X"FFFEFD",X"FFFEFF",X"FEFFFF",X"FCFFFF",X"FCFFFF",X"FEFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFCFF",X"FFFDFF",X"FFFFFF",X"FEFFFF",X"FCFFFD",X"FCFFFD",X"FEFFFD",X"FEFFFD",X"FEFFFB",X"FCFFFB",X"FCFFFD",X"FFFFFD",X"FFFBFF",X"FFF9FF",X"FFFDFF",X"F9FFFF",X"F4FFFF",X"FBFFFF",X"FFFFF8",X"FFFFFA",X"F8FFFF",X"F5FFFF",X"F8FFFF",X"FCFFFA",X"F1FFFF",X"F9FFFF",X"FFFDFF",X"FFFDFF",X"FCFFFF",X"F8FFFF",X"F9FFFF",X"FEFFFF",X"FFFFFB",X"FFFFFD",X"FFFEFF",X"FEFFFF",X"FCFFFF",X"FCFFFF",X"FFFFFF",X"FFFEFD",X"FEFFFF",X"FFFFFF",X"FFFFFB",X"FFFFFA",X"FFFFFB",X"FEFFFA",X"FEFFF4",X"FCFFF1",X"FEFEFF",X"FEFFFA",X"FEFFF3",X"FFFFF6",X"FFFFF8",X"FFFFF8",X"FFFFFD",X"FEFFFF",X"FFFDFF",X"FFFFFF",X"F9FFFB",X"F5FFFA",X"F5FFFA",X"F8FFFB",X"FCFFFF",X"FFFEFF",X"FBFFFF",X"FEFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFD",X"FFFFFD",X"FFFFFB",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFD",X"FEFFFD",X"F9FFFD",X"FBFFFD",X"FCFFFF",X"FEFFFF",X"FEFFFF",X"FCFFFF",X"FBFFFD",X"F9FFFD",X"FFFEFF",X"FFFFFF",X"FFFFFB",X"FFFFFB",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFF1",X"FFFFFF",X"FFFFFF",X"FFFFF4",X"FFFFF6",X"FFFDFF",X"FFFDFF",X"FFFFF6",X"FFFBFF",X"FFFEFF",X"FBFFFF",X"F8FFFF",X"F9FFFF",X"FCFFFF",X"FEFFFF",X"FFFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FCFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFD",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFDFF",X"FFFEFF",X"FFFEFF",X"FFFAFF",X"FFFEFF",X"F9FFFF",X"F9FFFF",X"FFFFFF",X"FFFEFF",X"FFFFFF",X"FBFFFF",X"FFFBFF",X"FFFAFF",X"FFFAFF",X"FFFEFD",X"F9FFFD",X"F8FFFD",X"FEFFFB",X"FFFDFB",X"F8FFFF",X"F9FFFF",X"FBFFFF",X"F9FFFF",X"F7FFFF",X"F7FFFF",X"F9FFFF",X"FCFFFF",X"FEFFFF",X"FEFFFF"),
(X"FEFFFF",X"FFFEFF",X"FFFDFF",X"FFF9FB",X"FFFEFF",X"FFFCFF",X"FCF0FC",X"FFF7FF",X"F7E3FE",X"E1D2E7",X"FEF8FF",X"FEFEFF",X"FEFFFD",X"FFFFFF",X"FFFDFF",X"FFFAFF",X"FFFFFD",X"FFFFFD",X"FCFBF9",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FFFEFF",X"FFFEFF",X"FEFEFE",X"FEFEFE",X"FFFFFF",X"FDFDFD",X"FFFFFF",X"F9F9F9",X"FFFFFD",X"FFFFFD",X"FBFFFB",X"FCFFFB",X"FEFFFF",X"FDFDFD",X"FBFBFB",X"FFFFFD",X"FDFFFA",X"FCFFFA",X"FFFBF6",X"FFFAF5",X"FFFFFB",X"F9FFFF",X"F7FFFF",X"F7FFFF",X"F8FFFF",X"F8FFFF",X"F8FFF8",X"FBFFFD",X"F9FFFD",X"FBFFFF",X"FCFFFF",X"FEFFFF",X"FBF9FE",X"FFFAFF",X"F8FFFF",X"FFFEFF",X"FFFBF8",X"FFFDFB",X"F7FAFF",X"F8FFFF",X"FCFFFF",X"FFFCF9",X"FCFCFA",X"FFFFFD",X"FBFDFC",X"FEFFFF",X"FEFFFF",X"FDFDFD",X"FDFCFA",X"FEFDF9",X"FBFFFA",X"FFFFFF",X"FEF9FF",X"FFFDFF",X"FCFFFB",X"FBFFFA",X"FDFDFD",X"FFFDFF",X"F8FFFB",X"FAFEFF",X"FBFAFF",X"FFFFFF",X"F9FEF8",X"FCFFF8",X"FFFFFB",X"FFFBFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"F8FEFE",X"F8FFFE",X"FCFFFD",X"FFFFFB",X"FFF8F6",X"FFFDFD",X"F8FEFC",X"F4FFFF",X"FFFAFD",X"FFF9FA",X"FFFFFD",X"FAFCF9",X"FBFBF9",X"FFFFFD",X"FBFFFA",X"F9FFFB",X"F8FFFF",X"FFFFFF",X"FFFDFF",X"FFFAFE",X"FDFDFF",X"FCFFFF",X"FBFCFE",X"FFFEFF",X"FBFFFE",X"FFFEFF",X"FFFEFF",X"FDFDFD",X"FBFFFF",X"F9FFFF",X"FCFFFF",X"FFFFFF",X"FDFDFD",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFDFF",X"FCFCFE",X"FEFFFF",X"FCFFFD",X"FAFBFD",X"FFFFFF",X"FBFBFB",X"FFFFFD",X"FFFFFD",X"FDFDFD",X"FBFBFB",X"FEFFFF",X"FCFFFF",X"FAFAF8",X"FFFFFA",X"FFFFFD",X"F6FAFD",X"FAFFFF",X"FEFFFF",X"FEF9FD",X"FFFDFF",X"FBFCFE",X"FAFFFF",X"FCFFFF",X"FCFAFD",X"FFFCFF",X"FFFFFF",X"FBFFFF",X"FFFDFF",X"FFFEFF",X"FBFAF8",X"FEFFFB",X"FBFFFA",X"FBFFFD",X"FAFFFE",X"FBFFFF",X"FDFFFA",X"F8FFFC",X"F7FFFD",X"FCFFFD",X"FCFBF9",X"FFFEFF",X"FFFFFF",X"FDFFFE",X"F8FFFF",X"FFFFFF",X"FFF9F6",X"FFFDFA",X"FFFEFF",X"F4F5F9",X"FEFFFF",X"FEFDFB",X"FFFFF3",X"FBF7F4",X"FFFCFF",X"FFFDFF",X"F5FAFE",X"F9FFFF",X"FBFFFF",X"FCFBFF",X"FEFFFB",X"FEFDF9",X"FFFDFD",X"FFFEFD",X"FFFFFD",X"FBFDFA",X"FFFFFD",X"FFFBFC",X"FDFFFC",X"FEFFFF",X"FFFEFF",X"FFFDFF",X"FFFCFF",X"FFFCFF",X"FCFBFF",X"FFFFFD",X"FCFFFF",X"F8FAF7",X"FEFFFA",X"FFFFFB",X"F9F9FB",X"FEFFFF",X"FCFFFF",X"F6FCFC",X"F8FCFD",X"FEFFFF",X"FFFFFD",X"FFFCF9",X"FFFEFB",X"FEFEFC",X"FBFDFC",X"FBFFFF",X"FCFFFF",X"FFFEFF",X"FFFDFF",X"FBF9FA",X"FBFFFD",X"F8FFFD",X"FAFFFE",X"FCFEFD",X"F5FFFF",X"FEFFFF",X"FFF9FF",X"FFF6FF",X"FFFDFF",X"FEFFFF",X"FEFFFD",X"FFFFFB",X"F7FCF8",X"FCFFFD",X"FEFFFF",X"FDFEFF",X"FAFBFD",X"FEFFFF",X"FCFFFD",X"FBFFFC",X"FFFCFF",X"FFFFFF",X"FFFFFB",X"FDFFFA",X"FDFDFF",X"FFFEFF",X"FFFEFD",X"FFFEFA",X"FBFFF1",X"F9FEFF",X"FCFEFF",X"FEFFFF",X"FEFFF7",X"FFFFFD",X"FFFEFF",X"FFFEFD",X"FEFCFF",X"FEFFFF",X"FAFBFD",X"FFFDFF",X"FFF6FC",X"FFFBFF",X"FEFCFF",X"FBFFFF",X"F9FFFF",X"FEFFFF",X"FFFBFC",X"FFFDFE",X"FEFEFE",X"FDFDFD",X"FFFDFF",X"FFFBFF",X"FFFFFF",X"FBFBFD",X"FFFEFF",X"FFFFFF",X"F7F7F9",X"FCFFFF",X"FBFFFF",X"F2FBF8",X"FFFEFF",X"FFFDFE",X"FFFEFF",X"FFFEFF",X"FCFCFC",X"FDFDFD",X"FFFFFF",X"FEFEFE",X"FEFFFA",X"FFFFFD",X"FFFDFF",X"FFF7FD",X"FFF7FD",X"FFFDFF",X"FFFEFF",X"FFFFFD",X"FFFDFF",X"F9F9FB",X"FEFFFF",X"FEFCFD",X"FFFCFD",X"FFFFFD",X"F5FBF7",X"F5FFFD",X"FCFFFF",X"FFFDFF",X"FFFDFF",X"FFFDFF",X"F4F4F6",X"FCFFFF",X"FCFEFD",X"FFFEFF",X"FFFEFF",X"FDF8FC",X"FFFDFF",X"FFFFFF",X"FCFFFF",X"FBFFFF",X"FEFFFF",X"FAF8F9",X"FDFFFE",X"FCFFFF"),
(X"F9FBFA",X"FFFEFF",X"FDF7F9",X"FFFDFF",X"FCFAFD",X"FFFDFF",X"F9EDF9",X"CDB8C9",X"523E59",X"44354A",X"F6F0FC",X"FEFEFF",X"F2F4F1",X"FFFFFF",X"FFFDFF",X"FFF8FF",X"F8F7F5",X"FEFDFB",X"FFFFFD",X"FEFDFB",X"FFFFFD",X"FBFAF8",X"FFFEFF",X"FFFDFE",X"FFFFFF",X"FDFDFD",X"FFFFFF",X"FDFDFD",X"FFFFFF",X"FBFBFB",X"FFFFFD",X"FEFEFC",X"FAFFFA",X"FAFFF9",X"FCFEFD",X"FDFDFD",X"FFFFFF",X"FFFFFD",X"FEFFFB",X"F9FEF7",X"FFF7F2",X"FFFDF8",X"FFFFFB",X"F8FFFE",X"F7FFFF",X"F7FFFF",X"F6FFFF",X"F9FFFF",X"FBFFFB",X"EFF5F1",X"FBFFFF",X"FBFFFF",X"F7FBFC",X"F6F7FB",X"FFFEFF",X"FFFDFF",X"F9FFFF",X"FFFBFC",X"FFF5F2",X"FFFAF8",X"FCFFFF",X"F7FFFF",X"FCFFFF",X"FFFDFA",X"FFFFFD",X"FFFFFD",X"FEFFFF",X"FDFEFF",X"FAFCFB",X"FEFEFE",X"FFFFFD",X"FFFFFB",X"FCFFFB",X"FCFCFE",X"FFFDFF",X"FEFCFF",X"FCFFFB",X"F5FCF4",X"FFFFFF",X"FFFDFF",X"F5FFF8",X"FCFFFF",X"FDFCFF",X"FFFFFF",X"FCFFFB",X"FAFFF6",X"F8F7F3",X"FFFCFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FBFFFF",X"F9FFFF",X"F8FDF9",X"FEFDF9",X"FFFDFB",X"FFFDFD",X"FBFFFF",X"EEFEFB",X"FFFAFD",X"FFFAFB",X"FEFDFB",X"FEFFFD",X"FFFFFD",X"FAFAF8",X"FBFFFA",X"F4FEF6",X"F9FFFF",X"FFFFFF",X"FFFAFE",X"FCF6FA",X"FFFFFF",X"FCFFFF",X"FBFCFE",X"FFFEFF",X"FBFFFE",X"FFFEFF",X"FCF8F9",X"FFFFFF",X"F4FAF8",X"F6FFFC",X"FCFFFF",X"F7F7F7",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"F8FDF9",X"FCFDFF",X"FCFCFC",X"FFFFFF",X"F9F8F6",X"FCFBF9",X"FFFFFF",X"FEFEFE",X"FEFFFF",X"FCFFFF",X"FAFAF8",X"FFFCF7",X"FEFDFB",X"F8FCFF",X"FBFFFF",X"FBFCFF",X"FFFDFF",X"FFFBFF",X"FCFDFF",X"FBFFFF",X"FCFFFF",X"FFFEFF",X"FFFDFF",X"FFFFFF",X"FAFEFF",X"FCF6FA",X"FFFEFF",X"FFFFFD",X"FEFFFB",X"FCFFFB",X"F5FBF7",X"FAFFFE",X"FBFFFF",X"FEFFFB",X"F8FFFC",X"F7FFFD",X"FBFFFC",X"FFFFFD",X"FFFEFF",X"FAFAFA",X"FDFFFE",X"F9FFFF",X"FFFFFF",X"FFFDFA",X"FFF8F5",X"FFFEFF",X"FEFFFF",X"FAFBFD",X"FFFEFC",X"FFFFF3",X"FFFEFB",X"FFFBFF",X"FAF8FF",X"FBFFFF",X"F9FFFF",X"FBFFFF",X"FFFEFF",X"FEFFFB",X"FFFFFB",X"FFFDFD",X"FAF6F5",X"FFFFFD",X"FCFEFB",X"FEFDFB",X"FFFCFD",X"F8FAF7",X"FEFFFF",X"FAF9FE",X"FEFBFF",X"FFFCFF",X"FFFCFF",X"FFFEFF",X"FFFFFD",X"FCFFFF",X"FEFFFD",X"FEFFFA",X"F9FAF5",X"FFFFFF",X"F7F8FD",X"F6FAFD",X"FBFFFF",X"FCFFFF",X"FCFEFD",X"FFFEFC",X"FDF9F6",X"FFFEFB",X"FFFFFD",X"FAFCFB",X"F6FCFC",X"FAFEFF",X"F6F4F5",X"FFFDFF",X"FFFEFF",X"F8FEFA",X"F2FDF7",X"FBFFFF",X"FEFFFF",X"F3FFFD",X"F5F6F8",X"FFFBFF",X"FFFAFF",X"FFFAFE",X"FEFFFF",X"F9FBF8",X"FFFFFB",X"FCFFFD",X"F9FEFA",X"FEFFFF",X"FAFBFD",X"FEFFFF",X"FEFFFF",X"F4F9F5",X"F9FEFA",X"FFFCFF",X"FDFDFD",X"FEFFFA",X"FEFFFB",X"FFFFFF",X"FFFDFF",X"FFFCFB",X"FFFCF8",X"FBFFF1",X"F4F9FC",X"FCFEFF",X"FAFCFB",X"FBFCF4",X"FFFFFD",X"FBF9FC",X"FFFEFD",X"FFFEFF",X"F8F9FB",X"F9FAFC",X"FFFDFF",X"FFFAFF",X"FFFCFF",X"FFFEFF",X"F6FCFC",X"F9FFFF",X"F6F8F7",X"FFFEFF",X"FFFEFF",X"FDFDFD",X"FFFFFF",X"FFFDFF",X"FFFAFE",X"FFFFFF",X"FFFFFF",X"FBF9FC",X"FFFFFF",X"FFFFFF",X"FBFFFF",X"FBFFFF",X"F8FFFE",X"FFFDFE",X"FCFAFB",X"FCFAFB",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFB",X"F7F6F4",X"FFFCFE",X"FFFBFF",X"FFFBFF",X"FAF4F8",X"FFFDFE",X"FCFCFA",X"FFFDFF",X"FFFFFF",X"F5F7F6",X"FDFBFC",X"FFFEFF",X"FAF9F7",X"FBFFFD",X"F3FFFB",X"F4F8F9",X"FBF9FC",X"FFFDFF",X"FFFDFF",X"FFFFFF",X"FAFEFF",X"F7F9F8",X"FFFEFF",X"FEFCFF",X"FFFDFF",X"FFFDFF",X"FCFCFE",X"F5F9F8",X"F6FCFA",X"FEFFFF",X"FFFEFF",X"FDFFFE",X"FCFFFF"),
(X"FFFFFF",X"F3F7F8",X"F6FCFC",X"FAF9FE",X"FFFBFF",X"E0CEDE",X"957E92",X"31192F",X"6D5877",X"BFB1B0",X"E1DCC8",X"FFFFF8",X"FFFEFF",X"FEFEFE",X"F9F8F6",X"FFFDFF",X"F5FFFA",X"F8FFFD",X"F7FBFC",X"FCFBFF",X"FDFCFF",X"FBFCFF",X"F7FCFF",X"F9FFFF",X"FAFAFA",X"FDFDFD",X"FFFEFF",X"F9F7F8",X"FFFDFF",X"FFFEFF",X"FFFDFF",X"FCF7FB",X"FBFDFA",X"F9FEFA",X"F9FEFA",X"FAFFFB",X"FBFDFA",X"FBFBFB",X"FEFAFB",X"FFF9FD",X"F2FFFF",X"F4FDFC",X"FFFAFF",X"FFF7FF",X"FFECFB",X"FFEFFF",X"FFF9FF",X"FFFBFF",X"FCF5FD",X"FFFDFF",X"FFFFFF",X"F7F9F8",X"F7F9F8",X"FFFFFF",X"FEFBFF",X"FAF4FF",X"FBFFFF",X"FFFDFD",X"FFF6EF",X"FFF8F1",X"FFFCFC",X"F7FAFF",X"FBFFFF",X"F4F8F9",X"FFFBF7",X"FBF7F4",X"FCFCFA",X"FEFFFF",X"F9FAFC",X"F9FBFA",X"FFFFFD",X"F2F1ED",X"F5FAF3",X"FFFAFF",X"FFF2FF",X"FFF8FF",X"FBF4FB",X"FBFBF9",X"F7F5F6",X"FFFBFF",X"F7F8FC",X"FFFBFF",X"FFF7FF",X"F8EEF9",X"FDFEF9",X"FCFFF6",X"FFFFFA",X"FFFBFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFBFF",X"FBF1F9",X"FFFAFF",X"FFFBFF",X"F9F4FB",X"FCF7FE",X"FFFBFF",X"FFF8FF",X"FFF0FC",X"FFFDFF",X"F5FFFF",X"F2F8F6",X"F9EFF0",X"FFF7FB",X"FFFCFB",X"FCFFFB",X"F7FDFD",X"FEFCFF",X"FFFCFF",X"FFFDFF",X"F6FCFC",X"F4FDFC",X"F8F9FB",X"FFF6FB",X"FFFEFF",X"FDF1F5",X"FFF3FA",X"FFF9FF",X"F9F5F6",X"FAFFFE",X"FAFFFE",X"FEFFFF",X"FDFEFF",X"F9F9FB",X"FBF9FA",X"FAF8F9",X"FBF9FA",X"FEFFFF",X"FBFEFF",X"F3FAFF",X"FEFFFF",X"F6F6F8",X"FFFDFC",X"FFFEFB",X"FFFBF8",X"FFFEFD",X"FDFDFF",X"FBFCFF",X"F6FBFE",X"FFFCF6",X"FFFDEF",X"FFF9ED",X"FFFEFA",X"FAF9FE",X"F9F6FF",X"FFFBFF",X"FAF4F8",X"FAFBFD",X"FAFFFF",X"FCFDFF",X"FFFAFE",X"FFFAFE",X"F5FEFD",X"EBFFFB",X"F2FFFF",X"F6FFFF",X"F7FBFA",X"F9F5F4",X"FAEFF3",X"FFFAFF",X"FFF9FF",X"FFF3FF",X"FFF1FE",X"FFF7FF",X"FFFAFF",X"F6F4F9",X"FBFFFF",X"F4FFFF",X"F3FEFA",X"FEF8FA",X"F5F9FC",X"F6F9FE",X"FFFEFF",X"FFFAFE",X"FFF7FA",X"FFFDFF",X"F7F8FC",X"F7FFFF",X"FFF9F6",X"FFFDFF",X"F3F9FF",X"EFFCFF",X"F8FFFF",X"FCFDFF",X"F9F6FD",X"FFFBFF",X"EBFBFB",X"F6FAFB",X"FFFCFD",X"FFF9F8",X"FFFFFA",X"FAFCF7",X"FBFBFB",X"FFFBFF",X"FCFFFD",X"FFFFFA",X"F4F4EC",X"FFFEFA",X"FEF6F4",X"F3EBE9",X"FFFFF6",X"FEFAEE",X"F8F9EB",X"F9F8F4",X"FFFBF8",X"FFFEF5",X"FFFEFF",X"F9F7FF",X"FCFFFF",X"FAFFEC",X"FBFFFF",X"FAFAFC",X"FFFAFF",X"FFF5FE",X"FFF2FC",X"FFF9FF",X"F8F6F9",X"FEFFFF",X"FEFFFF",X"FDF9FA",X"FFFDFF",X"F5F5F5",X"F4FFFB",X"F7FFFF",X"FBFCFF",X"FFFBFF",X"F9FFFF",X"F7F8FC",X"FCFBFF",X"FFFEFF",X"F5F6FA",X"FCFFFF",X"FCFCFA",X"FFFEFB",X"FFF6F7",X"FFFDFF",X"FAF5F9",X"FEFDFF",X"FCFBFF",X"FFFCFF",X"FEF8FA",X"FFFCFD",X"FFFDFF",X"FEFCFD",X"FDFEF9",X"FEFFFF",X"FFFEFF",X"FCFAFB",X"FFFDF2",X"FFFFEA",X"FFFFF3",X"FEFEF6",X"FFFFFD",X"FFFEFF",X"FFFEFF",X"FDFCF7",X"F5F4F0",X"FCFAFB",X"F2FCFB",X"F2FFFE",X"F7FFFF",X"F4F8F9",X"F8F2F6",X"FFFCFF",X"FFFFFF",X"F8FFFF",X"F4FDFA",X"FFFFFF",X"FFF9FB",X"FEFAFB",X"FBFFFE",X"F2F8F6",X"F6F4F5",X"FFFBFF",X"FDF7FB",X"FFFCFF",X"FFF6FA",X"FFF9FD",X"FFFAFE",X"FAF1F4",X"FBF5F5",X"FFFBFA",X"FFFCFD",X"FFFEFF",X"FFFDFE",X"FAF8F9",X"FCFAFB",X"FEFEFE",X"FDFDFD",X"FDFDFD",X"F9FAFC",X"FEFFFF",X"F8FCFD",X"FAFEFD",X"FAFEFD",X"FCFFFF",X"FEFFFD",X"F7F9F6",X"F2F8F8",X"FFFFFF",X"FFFDFF",X"FDF4F7",X"FFFEFD",X"FFFFFD",X"F8F4F1",X"FFFEFB",X"F5FFFF",X"F7FFFF",X"F3F9F9",X"FFFCFF",X"FFFBFF",X"FDF8FE",X"FBFFFF",X"EFFFFE",X"FAF9FE",X"FEFCFF",X"FFFAFF",X"FFFEFF",X"FEFFFF",X"FFFFFF",X"FFF9FB",X"FFF7FB",X"FEF5F8",X"FFFAFC"),
(X"FDFDFF",X"F7FBFC",X"FAFFFF",X"FCFBFF",X"FFF5FE",X"BBA9B9",X"DCC5D9",X"FCE4FA",X"FEE9FF",X"FBEDEC",X"FFFFEC",X"FFFEF7",X"FAF8FD",X"FFFFFF",X"FEFDFB",X"FFFDFF",X"EFFFF4",X"F6FFFB",X"F8FCFD",X"F8F7FD",X"FFFEFF",X"FEFFFF",X"F5FAFD",X"F9FFFF",X"FDFDFD",X"FAFAFA",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FCFAFD",X"FAF5F9",X"FDF8FC",X"FCFEFB",X"FAFFFB",X"FAFFFB",X"FCFFFD",X"FEFFFD",X"F8F8F8",X"FFFBFC",X"FFFDFF",X"F1FFFE",X"F6FFFE",X"FEF5FA",X"FFF7FF",X"FFF3FF",X"FFF6FF",X"FFF7FF",X"F4EDFD",X"FFFCFF",X"FEF9FF",X"FCFCFE",X"FEFFFF",X"F9FBFA",X"FEFEFF",X"FFFDFF",X"FFFCFF",X"F5FAFF",X"FFFDFD",X"FFF3EC",X"FFFBF4",X"FEF8F8",X"F3F6FB",X"F9FEFF",X"FCFFFF",X"FFFEFA",X"FFFBF8",X"F7F7F5",X"FCFDFF",X"FCFDFF",X"FBFDFC",X"FFFFFD",X"FFFFFB",X"FCFFFA",X"FFFBFF",X"FFF3FF",X"FCEBFD",X"FFFCFF",X"FFFFFD",X"FFFEFF",X"FFFAFF",X"FEFFFF",X"FDF5FF",X"FFF7FF",X"FFF8FF",X"FFFFFB",X"F8FEF2",X"FCFBF6",X"FFF6FA",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFCFF",X"F8EEF6",X"FFFAFF",X"FFFAFF",X"FFFBFF",X"FFFDFF",X"F6ECF4",X"FFF5FE",X"FFF6FF",X"FAF5FB",X"F7FFFF",X"FBFFFF",X"FFFCFD",X"FFF8FC",X"FCF2F1",X"F9FEF8",X"FBFFFF",X"F6F4F7",X"FFF7FC",X"FFFDFF",X"F4FAFA",X"F6FFFE",X"FEFFFF",X"FFF7FC",X"FFFEFF",X"FEF2F6",X"FFF8FF",X"FFF9FF",X"FFFEFF",X"F7FDFB",X"F4FAF8",X"F7F9F8",X"FBFCFF",X"FAFAFC",X"FFFEFF",X"FFFDFE",X"FAF8F9",X"FCFDFF",X"FCFFFF",X"F8FFFF",X"FBFCFF",X"FFFFFF",X"FDF9F8",X"FFFAF7",X"FAF5F2",X"FDF9F8",X"FFFFFF",X"FAFBFF",X"F7FCFF",X"FDF8F2",X"FFFDEF",X"FFFAEE",X"FFFAF6",X"FDFCFF",X"F7F4FD",X"FFFBFF",X"FFFCFF",X"FEFFFF",X"FBFFFF",X"FEFFFF",X"FFFBFF",X"FFFBFF",X"F7FFFF",X"EFFFFF",X"EFFFFE",X"F4FFFE",X"FAFEFD",X"FFFEFD",X"FFFAFE",X"FFF2F9",X"FFF0FB",X"FFF6FF",X"FFF7FF",X"FFFAFF",X"FFFCFF",X"FFFDFF",X"F7FDFD",X"ECFDF7",X"F4FFFB",X"FFFDFF",X"FCFFFF",X"F7FAFF",X"FBFAFF",X"FFFDFF",X"FFFAFD",X"FDF7F9",X"FEFFFF",X"F6FFFF",X"FFF6F3",X"FDF8FC",X"F7FDFF",X"F5FFFF",X"F8FFFF",X"FBFCFF",X"FDFAFF",X"FFFBFF",X"F4FFFF",X"F9FDFE",X"FFFCFD",X"FFFBFA",X"F8F7F2",X"FAFCF7",X"FFFFFF",X"FFFBFF",X"F5FAF6",X"F6F7F1",X"FFFFF8",X"FFFAF6",X"FCF4F2",X"FFFDFB",X"FFFFF6",X"FFFDF1",X"FFFFF3",X"FCFBF7",X"FFFCF9",X"FFFDF4",X"FCFAFB",X"FBF9FF",X"FAFEFF",X"F2FCE4",X"F4FAFA",X"F8F8FA",X"FFF7FF",X"FFFAFF",X"FFF9FF",X"FFFBFF",X"FBF9FC",X"F8F9FB",X"FBFCFE",X"FFFDFE",X"FEF8FA",X"FEFEFE",X"F8FFFF",X"F7FFFF",X"F5F6FA",X"FFFBFF",X"F1FAF9",X"FEFFFF",X"F7F6FC",X"FFFEFF",X"FAFBFF",X"FCFFFF",X"FDFDFB",X"FAF6F3",X"FFFCFD",X"FDF7F9",X"FCF7FB",X"FDFCFF",X"FFFEFF",X"F5F0F4",X"FFFDFF",X"FFF7F8",X"FFFCFF",X"FFFDFE",X"FFFFFB",X"FEFFFF",X"FDFCFF",X"FBF9FA",X"FEFAEF",X"FFFEE8",X"F7F7EB",X"FFFFF8",X"F4F3F1",X"FFFDFF",X"FFFEFF",X"FAF9F4",X"FFFEFA",X"FFFEFF",X"F7FFFF",X"F5FFFF",X"E7F3F1",X"F9FDFE",X"FFFDFF",X"F9F0F5",X"FCFCFE",X"F5FFFE",X"F3FCF9",X"FFFFFF",X"FFFDFF",X"FEFAFB",X"F2F6F5",X"FBFFFF",X"FFFEFF",X"FDF2F6",X"FDF7FB",X"FFF8FD",X"FFF8FC",X"FFF6FA",X"FFFAFE",X"FFFCFF",X"FFFCFC",X"FFFEFD",X"FCF8F9",X"FFFCFD",X"FFFBFC",X"FEFCFD",X"FFFEFF",X"FEFEFE",X"FAFAFA",X"FCFCFC",X"FCFDFF",X"FCFDFF",X"FCFFFF",X"F5F9F8",X"FCFFFF",X"F7FBFA",X"F2F4F1",X"FEFFFD",X"FBFFFF",X"FEFEFF",X"FBF5F7",X"FFFAFD",X"FFFEFD",X"FEFDFB",X"FEFAF7",X"FFFEFB",X"EAF9F6",X"F7FFFF",X"F8FEFE",X"FFFDFF",X"FDF3FB",X"FEF9FF",X"F6FBFE",X"F2FFFF",X"FFFEFF",X"FFFEFF",X"FAF5FB",X"FDFBFE",X"F9FAFC",X"F2F2F2",X"FFFBFD",X"FFF8FC",X"FFFCFF",X"FDF7F9"),
(X"FAFBFD",X"F4FFFF",X"EEFFFF",X"EAF5F7",X"FFF2FF",X"FFEDFF",X"FFE8FF",X"FFF5FF",X"FFF8FF",X"FFFFD4",X"FFFFB9",X"FFFBE1",X"FFFCFF",X"FFFCFB",X"F9FAF2",X"FEFFFF",X"F7FFFA",X"F7F9F8",X"FFFAFF",X"FFEEFF",X"FFF3FF",X"FFF1FF",X"FFF7FF",X"F9F6FF",X"FFFFFD",X"FAF9F7",X"F7F5F6",X"FAF5F9",X"FEF9FF",X"FFFCFF",X"FEF7FF",X"FFFBFF",X"FFFCFF",X"FFFEFF",X"F9FBFA",X"FCFFFD",X"FFFFFF",X"FFF5FE",X"FFF4FF",X"FFEFFF",X"F8F1FF",X"FFF6FF",X"FFE5FF",X"FFDFFF",X"FFD2F6",X"FFD6FC",X"FFE0FF",X"FFEAFF",X"FFE1FF",X"FFF2FF",X"FFEEFE",X"FBEFF1",X"FFFFFA",X"FFFFFB",X"FDFDFD",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFF9F2",X"FFF0D8",X"FFF1C6",X"FFE8B4",X"FFEDC0",X"FFEDCA",X"F8EDE7",X"FFFEF8",X"FFFEFB",X"FDFDFD",X"FEFFFF",X"F7F8FA",X"F8F8F8",X"FEFDFB",X"FAFBF6",X"FFF1FF",X"FFE3FF",X"FFE5FF",X"FFEAFF",X"F7E9F6",X"F5E7F4",X"FFF4FF",X"FFEAFF",X"FFDFFF",X"FFE3FF",X"FFEDFF",X"FFFCFF",X"FAFFF6",X"FEFFFB",X"FFFBFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFE3F8",X"FFE5FF",X"FFD6FF",X"FFC1F2",X"FFDAFF",X"FFD5F9",X"FFDFFE",X"FFE0FD",X"FFE9FF",X"FFE9FF",X"FFF2FF",X"FFF1FE",X"FFFEFF",X"F1FAF9",X"FBFFFF",X"F9FEFA",X"FEFFFF",X"FEF9FD",X"FFF8FD",X"FFFFFF",X"F7FFFF",X"F6FFFF",X"F7F7F9",X"FFF9FF",X"FDECF2",X"FFF0FB",X"FFE1EF",X"FFE4F1",X"FFEFF6",X"FFFEFF",X"FEFFFF",X"FCFCFC",X"FBFEFF",X"FBFCFF",X"FBFBF9",X"FFFEFA",X"FAFAF8",X"FBFFFF",X"F9FFFF",X"ECF3FF",X"F9F8FD",X"FEFCFF",X"FAF4F4",X"FAF2F0",X"FFFDFB",X"FEF8F8",X"FCFAFD",X"FAF9FE",X"FBFDF8",X"FFF3E3",X"FFF2D7",X"FFF5DA",X"FFF1E3",X"FDF3F2",X"FFFBFF",X"FFF7FF",X"FAF4F8",X"F8F8FA",X"F8FCFD",X"FFFDFF",X"FFFCFF",X"FFFEFF",X"F1FFFF",X"D9FFF4",X"CDFFFB",X"D7FFFB",X"EAFCFC",X"FFFAFF",X"FFE5F9",X"FFE1FF",X"FFDBFF",X"FFD3FE",X"FFD4FD",X"FFDAFF",X"FFD0FA",X"FFDAFF",X"FFE5FE",X"F9F6FD",X"F8FFFF",X"F6F1F5",X"E9FFFF",X"DBFEFF",X"D9FFFF",X"E5FFFF",X"F0FFFC",X"EDFCF5",X"E8FFFF",X"D0FFFF",X"C2FFFF",X"B8FFFF",X"BEFFFF",X"C6FFFF",X"D1FAFF",X"D6FBFF",X"CBFEFF",X"C7FFFF",X"DBFCFF",X"F3FFFF",X"FEF9FF",X"FFFAFB",X"FFFEFA",X"F7FDFB",X"F4F9FD",X"F5F5FF",X"F3F5FF",X"FFFFF6",X"FFFFDA",X"FFFFBC",X"FFFFB1",X"FFFFA5",X"FEFFA2",X"FFFFA6",X"FFFFAF",X"FFFFC2",X"FFFCBA",X"FFFFAD",X"FFFFCB",X"FFFBFF",X"F9F5FF",X"FBFCFE",X"FBF9FA",X"FFFBFF",X"FCF0FE",X"FEEDFF",X"FFF6FF",X"F8E6F6",X"FFF9FF",X"FFF7FB",X"F4F8F7",X"FFFEFF",X"FBF5F7",X"FFFFFF",X"EBF4F3",X"F2F3F7",X"FFF6FF",X"FFE4FC",X"FFF0FD",X"FBFFFF",X"E7FFFF",X"D3FAF5",X"F1FFFF",X"FFFEFF",X"FFFCFE",X"FFFFFB",X"FBF5F5",X"FAFAFC",X"F9FFFF",X"EFFDFE",X"F2FFFF",X"F9FFFF",X"F6F6F8",X"FBF5F5",X"FFFDFF",X"FFFFFD",X"FBFCF7",X"F7F8FA",X"FEFDFF",X"FFFEFD",X"FFFFEA",X"FEFBD0",X"FFFFCD",X"FFFFB3",X"FFFCB1",X"FFFFDE",X"FFF8F9",X"FEFDFB",X"F5F7F2",X"FAFEFF",X"F1FBFA",X"D9FFF7",X"BEFFF2",X"B9FFF6",X"B7FFE9",X"E3FFFF",X"EFFEFB",X"FCFDFF",X"FCFFFF",X"F8F4F5",X"FFF9FC",X"FEFCFD",X"F5FFFF",X"F0FFFF",X"EAFBF5",X"F7FFFD",X"FFFBFF",X"FBEAF0",X"FFF2FA",X"FFE6EE",X"FFDBE5",X"FFE7EF",X"FFE7EF",X"FFEFF6",X"FFFBFD",X"FFFAFC",X"FFFBFC",X"FFFDFE",X"FFFDFE",X"FAFAFA",X"FAFAFA",X"FEFFFF",X"FEFCFF",X"EFF8FF",X"E1FAFF",X"D9FCFF",X"D9FCFF",X"E3FDFF",X"F6FFFF",X"F9F8F3",X"F8FFFF",X"F6F4F7",X"FFFAFD",X"FFFEFF",X"F3F5F2",X"FFFEFB",X"FFE9F0",X"FFD6E6",X"FFE4F3",X"FFE1E9",X"FFFAF9",X"F7F7F5",X"FFFEFF",X"FFFDFF",X"F2FAFC",X"F0FFFF",X"D4F9F2",X"E3FFFE",X"E9FFFF",X"E6FFF9",X"F1FFFF",X"F7FFFF",X"F6F6F6",X"FFFAFB",X"FFE6F1",X"FFF6FF"),
(X"E8E9EB",X"9FAFAE",X"5F7874",X"5F6A6C",X"726473",X"7E5E76",X"765874",X"594560",X"554353",X"A29B6D",X"D1D18B",X"E5DFC5",X"FFFCFF",X"F9F5F4",X"FFFFF8",X"FBFCFF",X"F5FFF8",X"FAFCFB",X"FBEFFD",X"FFF2FF",X"F6DBFA",X"C2AEC9",X"695E6F",X"585560",X"3C3B39",X"302F2D",X"464445",X"645F63",X"635E64",X"645D65",X"7D767E",X"BAB2BD",X"F3ECF4",X"FFFEFF",X"FAFCFB",X"F7FCF8",X"FAFAFA",X"FFF9FF",X"FFF7FF",X"FFEAFF",X"EAE3FF",X"B4A3C5",X"846587",X"7B4E6F",X"4D193D",X"4F1D43",X"754B73",X"88628B",X"B892BB",X"F6D7F6",X"FFF0FF",X"FFFBFD",X"FFFCF7",X"FFFFFB",X"FAFAFA",X"FFFEFF",X"FFFEFF",X"F9F7F8",X"DED5CE",X"A98B73",X"BE8D62",X"CA9561",X"D2A77A",X"B79D7A",X"C0B5AF",X"F4EDE7",X"FFFCF9",X"F9F9F9",X"FEFFFF",X"FEFFFF",X"FDFDFD",X"FFFFFD",X"FBFCF7",X"A08DA0",X"6C466F",X"916B94",X"7E647F",X"817380",X"6F616E",X"665366",X"7E6481",X"8E6A90",X"805985",X"A98FAC",X"FFFAFE",X"FBFFF7",X"F8FAF5",X"FFFCFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"C3A3B8",X"854E6E",X"B56693",X"B96798",X"B3709C",X"996589",X"905D7C",X"9F6784",X"B18DA7",X"EBC9E1",X"F8DDF0",X"FFF9FF",X"F9F8FD",X"F1FAF9",X"FBFFFF",X"F7FCF8",X"F5F6F8",X"FFFDFF",X"FFFCFF",X"F3F3F5",X"EBF7F5",X"AAB6B4",X"59595B",X"5D4E55",X"604F55",X"5D3D48",X"805664",X"8B6572",X"826D74",X"CDC9CA",X"ECEEED",X"FFFFFF",X"F9FCFF",X"FEFFFF",X"F7F7F5",X"FFFFFB",X"FFFFFD",X"EEF2F5",X"C0C7D1",X"6F7686",X"616065",X"666467",X"6C6666",X"847C7A",X"D5CDCB",X"FFF9F9",X"FFFEFF",X"F9F8FD",X"F1F3EE",X"CDC1B1",X"B3997E",X"CEB398",X"B7A597",X"514746",X"C9BEC6",X"FFF3FD",X"FFFDFF",X"FFFFFF",X"FCFFFF",X"FFFDFF",X"FFF9FE",X"F7F5F8",X"C0D3CF",X"7BA196",X"67A195",X"79A49D",X"758787",X"C8BCC6",X"866377",X"9A6484",X"A6688F",X"A4638E",X"A56891",X"A3628A",X"A45781",X"B4688F",X"91657E",X"5D5A61",X"5F696A",X"6A6569",X"7C9693",X"83A6AC",X"789EAB",X"B7D4DC",X"F5FFFF",X"F5FFFD",X"A1BFC1",X"6E9EAA",X"6FB1C9",X"58A2BB",X"61ACC1",X"71ACBA",X"6F989E",X"779CA2",X"72A5B6",X"5295AF",X"A2C3CC",X"F3FFFF",X"FEF9FF",X"FFF6F7",X"FFFFFB",X"F6FCFA",X"F3F8FC",X"FEFEFF",X"FAFCFF",X"E1E3D8",X"DFE2B7",X"D2D38F",X"DAD986",X"D3D379",X"D0D174",X"CACE70",X"D1D080",X"D0CC8F",X"D8D391",X"E2E18E",X"D3D09B",X"DDD5E0",X"FFFBFF",X"FEFFFF",X"FFFEFF",X"878087",X"584C5A",X"79687A",X"6D5A6D",X"7B6979",X"65555F",X"E5D9DD",X"FCFFFF",X"F1EFF0",X"FFFDFF",X"FDFDFD",X"F9FFFF",X"EAEBEF",X"796473",X"815971",X"775F6C",X"565B5F",X"6A8D89",X"739A95",X"D6EAEB",X"F8F7FC",X"FCF6F8",X"FFFFFB",X"FAF4F4",X"FFFFFF",X"8F9799",X"8D9B9C",X"F1FFFF",X"F3FBFD",X"F7F7F9",X"FFFDFD",X"FDF8FE",X"FEFDFB",X"FFFFFB",X"FEFFFF",X"FFFEFF",X"F8F4F3",X"D4CFB9",X"AFAC81",X"C0AE7C",X"C8BD6E",X"C8C075",X"9D9473",X"A69D9E",X"FDFCFA",X"FEFFFB",X"F4F8F9",X"E0EAE9",X"729C90",X"76C1AA",X"5DB69A",X"6CB49E",X"729C90",X"C7D6D3",X"FBFCFE",X"F4F8F7",X"FFFEFF",X"FDF4F7",X"FFFEFF",X"EDFCF7",X"E3FAF2",X"F4FFFF",X"E1EAE7",X"A4989C",X"76656B",X"6D565E",X"684951",X"6B4751",X"815C64",X"856068",X"88656C",X"D1CBCD",X"E7E1E3",X"FDF9FA",X"FEFCFD",X"FAF8F9",X"FFFFFF",X"FFFFFF",X"F8FAF9",X"DBD9DE",X"6C7584",X"607998",X"6386B0",X"6184AC",X"516B84",X"B1BCC2",X"FAF9F4",X"F7FFFF",X"FFFEFF",X"FFF6F9",X"FDF9FA",X"FEFFFD",X"DED9D6",X"89666D",X"A46777",X"A16372",X"87626A",X"716766",X"F1F1EF",X"FCF8F9",X"FCF7FB",X"D6DEE0",X"677B79",X"84A9A2",X"81A19C",X"76918C",X"68817B",X"4D625D",X"47534F",X"646464",X"6D6465",X"7E5E69",X"EFD4DD"),
(X"FBFFFF",X"C6E1DC",X"234B43",X"000607",X"08000B",X"482440",X"B091B0",X"8B7B96",X"211310",X"9C9B49",X"BBBE53",X"FFFED2",X"FFF7FD",X"FFFEF9",X"FBFDEF",X"F5F8FD",X"FFFBF7",X"FFF8FF",X"FFE9FF",X"D39DCE",X"480D43",X"3D0939",X"5C3759",X"8C7089",X"B6B2B1",X"C5C1C0",X"AEAAAB",X"585357",X"0B040C",X"040007",X"060009",X"08000B",X"E2D1E4",X"FFF6FF",X"FFFEFF",X"F9FBFA",X"FFFEFF",X"FFF8FF",X"FBDCFB",X"C79EC6",X"740060",X"56004D",X"5E2260",X"AF93BC",X"D0C1E2",X"D9BFE6",X"A678A9",X"51144F",X"49084A",X"460D40",X"9D7492",X"ECD5DB",X"FEF5EE",X"FFFFF6",X"FDFFF9",X"FBFFFC",X"FDFAF3",X"FBFFFF",X"F7F4EB",X"D7A87C",X"E48126",X"F17503",X"E0770E",X"D38532",X"E8DBD2",X"FFFCF6",X"FFFEFB",X"F8F8F8",X"F8F9FD",X"F9FAFE",X"FBFBFD",X"FCFAFB",X"FEFAF9",X"EAD0EB",X"B481B9",X"3F0744",X"380F39",X"10000F",X"5B455A",X"B096AF",X"855181",X"4D124C",X"3A003C",X"9D749E",X"FFF3FF",X"F6FBF5",X"FCFFFF",X"FCF9FF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"EDD5ED",X"DA82B5",X"AC065C",X"CB076B",X"AF025E",X"C84F96",X"EB9CCC",X"94567B",X"8C0347",X"B10F5B",X"E33F88",X"FFAEE1",X"FFF3FF",X"F3FFFF",X"F6FBFE",X"FFF7FF",X"FDFDFF",X"FFF9FD",X"F3EDF1",X"B3B7B8",X"596966",X"000805",X"010002",X"907C85",X"C9AEB7",X"DFB3C2",X"C08599",X"531C2F",X"160000",X"080000",X"3B393A",X"D1CFD0",X"F1F3FF",X"FEFFFF",X"F4F4F2",X"FAFAF2",X"FFFFFB",X"FCFFFF",X"E2EAF7",X"7E869D",X"060409",X"030002",X"060000",X"B5ABAA",X"FFF9F8",X"FFFBFC",X"F5F0F4",X"FFFEFF",X"FCFCF2",X"FFF0D8",X"DBB892",X"AF8763",X"4B2F19",X"130000",X"9A878B",X"FFF6FD",X"FEF8FC",X"FBFBFD",X"FDFEFF",X"FFFAFE",X"FFFBFF",X"FFFFFF",X"A3BCB6",X"245446",X"48A392",X"1E6257",X"9BB7BA",X"A493A5",X"270012",X"711D4F",X"720C4B",X"871A5E",X"78205D",X"88165B",X"A50A58",X"AE0755",X"7D083F",X"1F0011",X"000007",X"0D0C12",X"05080F",X"00081F",X"011A39",X"BDC9E1",X"F8EEF7",X"FFFBFD",X"ECF5FF",X"94B5D6",X"0083C1",X"23A8E1",X"2291BF",X"569CBE",X"96BED7",X"7CAAC4",X"3C96B9",X"078AB6",X"89B7C7",X"EDFFFF",X"FDFBFF",X"FDF4F7",X"FBFBF9",X"F4FEFD",X"F7FFFF",X"ECF3FF",X"A9ACB3",X"000300",X"979B5E",X"E4E78C",X"CDCD6B",X"E4DF8D",X"ECE4A5",X"EBE3B2",X"E2DC7A",X"D3C972",X"D0CB53",X"D0D62E",X"9A9D18",X"8D8763",X"FFF8FF",X"FBFAF5",X"FBFFFE",X"E6BCD0",X"C96192",X"920040",X"A1074D",X"67002A",X"C490A7",X"FFF7FA",X"F9FFFD",X"FFFFFF",X"FFFEFF",X"FFFFFF",X"F3F4F6",X"FFF6FF",X"DEB6CE",X"4A0A2D",X"2E0010",X"000205",X"074B3C",X"65B2A2",X"DDFFFC",X"FFFDFF",X"FFF9FD",X"F8F9F4",X"F9FFFF",X"E7F7F4",X"64817D",X"000B07",X"799D99",X"E4FFFD",X"F4FFFF",X"F3FCF9",X"FFFDFF",X"FFFFFD",X"FBFBF9",X"F9FAFE",X"FEFDFF",X"FFFBF8",X"F2EFD0",X"E1DEA7",X"CFB044",X"AD9B00",X"B7AD0D",X"D6CB7B",X"E0D6CD",X"FFFEFF",X"F4FAF6",X"F8FFFF",X"F1F5F6",X"96DAC5",X"0CA070",X"07C587",X"00A972",X"63CCAB",X"DCFDF4",X"FFFBFF",X"FEFEFE",X"FFFCFF",X"FBF0F4",X"FEFFFF",X"ECFFFB",X"E2FFFB",X"AECFC4",X"000900",X"0D0002",X"553E46",X"B5949D",X"ECBECB",X"DFA9B7",X"AE7181",X"733343",X"440414",X"040000",X"3F393B",X"AEAAAB",X"FCF8F9",X"FFFEFF",X"F6F6F6",X"FBFBFB",X"FEFFFF",X"FBF5F9",X"AEBBDD",X"00105D",X"124DB5",X"00379D",X"5981C6",X"E3F2FF",X"FFFFF4",X"EDF7F6",X"FFFEFF",X"FFF9FC",X"FCFEFD",X"F2FDF7",X"FFF7F6",X"ECADBE",X"700523",X"A50026",X"73001D",X"DDB6BB",X"F8FDF6",X"F9FFFB",X"FBFDFC",X"F2F6F7",X"B9C5C3",X"3A5350",X"000505",X"000304",X"0C0D11",X"5E555A",X"6F5860",X"200005",X"420F1E",X"431021",X"F7C8D8"),
(X"F9FEFF",X"E8FFFE",X"608880",X"000607",X"0B000E",X"C7A3BF",X"FFE9FF",X"FFF6FF",X"FEF0ED",X"EFEE9C",X"BFC257",X"EFE8BC",X"FFFBFF",X"FCF9F4",X"FDFFF1",X"FCFFFF",X"FFFAF6",X"FCEBF5",X"A47D9C",X"380233",X"A0659B",X"FAC6F6",X"FFE4FF",X"FFF0FF",X"FFFEFD",X"FCF8F7",X"FFFBFC",X"FEF9FD",X"EDE6EE",X"C5BDC8",X"5A4F5D",X"130816",X"E1D0E3",X"FFF9FF",X"FFFDFF",X"F6F8F7",X"FFFEFF",X"F7E6F6",X"A98AA9",X"330A32",X"80086C",X"F797EE",X"FFD4FF",X"FFE8FF",X"FEEFFF",X"FFF3FF",X"FFE4FF",X"FFD2FF",X"C685C7",X"3C0336",X"1B0010",X"20090F",X"EBE2DB",X"FFFFF5",X"F7FAF3",X"FCFFFD",X"FEFBF4",X"F9FFFF",X"FDFAF1",X"FFE5B9",X"F8953A",X"F07402",X"E0770E",X"FFD481",X"FFF7EE",X"FFFCF6",X"FFFBF8",X"FEFEFE",X"FEFFFF",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFDFC",X"FFEEFF",X"FDCAFF",X"35003A",X"1A001B",X"40263F",X"ECD6EB",X"FFEDFF",X"FFE1FF",X"FFC5FF",X"824684",X"855C86",X"FFF8FF",X"FCFFFB",X"F6FAF9",X"FFFDFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFF4FF",X"FFBEF1",X"B50F65",X"DD197D",X"BD106C",X"FF9AE1",X"FFDDFF",X"FFD8FD",X"FF83C7",X"A80652",X"B10D56",X"AE3F72",X"FFE0F5",X"F4FFFF",X"FAFFFF",X"FFF4FE",X"FFFFFF",X"F3EDF1",X"938D91",X"000102",X"0D1D1A",X"AFBEBB",X"F5F3F6",X"FFEFF8",X"FFF5FE",X"FFEDFC",X"FFE1F5",X"FFD1E4",X"B5949F",X"0A0002",X"050304",X"010000",X"BBBDC9",X"FBFCFF",X"FFFFFD",X"FFFFF8",X"F6F7F2",X"FAFDFF",X"F8FFFF",X"9FA7BE",X"010004",X"2D282C",X"0D0405",X"EFE5E4",X"FEF4F3",X"FFFCFD",X"FFFDFF",X"FDFBFF",X"FEFEF4",X"FFF8E0",X"FFF0CA",X"E0B894",X"160000",X"321F19",X"251216",X"F5E0E7",X"FFFCFF",X"FEFEFF",X"FEFFFF",X"FCF7FB",X"FFFAFF",X"FFFFFF",X"88A19B",X"001103",X"328D7C",X"A4E8DD",X"E9FFFF",X"4F3E50",X"9A6285",X"FEAADC",X"FFC4FF",X"FFBEFF",X"FFCAFF",X"FFC3FF",X"FF6CBA",X"AC0553",X"C24D84",X"FFDDF7",X"F6F6FE",X"E6E5EB",X"D0D3DA",X"96A6BD",X"000524",X"AAB6CE",X"FFFBFF",X"FFF7F9",X"F3FCFF",X"BBDCFD",X"0690CE",X"169BD4",X"48B7E5",X"BBFFFF",X"DDFFFF",X"CFFDFF",X"ACFFFF",X"22A5D1",X"8AB8C8",X"E5FCFF",X"F9F7FF",X"FFFCFF",X"FBFBF9",X"F7FFFF",X"E8F2FB",X"949BAD",X"000007",X"010400",X"C5C98C",X"FFFFA9",X"FFFFA1",X"FFFFAE",X"FFFFC3",X"FFFFCE",X"FFFFA1",X"FFFFAC",X"FDF880",X"F2F850",X"AFB22D",X"716B47",X"FEF6FF",X"FFFFFA",X"F7FBFA",X"FFF0FF",X"FFAADB",X"A10A4F",X"C3296F",X"A43367",X"FFD3EA",X"FFFCFF",X"FAFFFE",X"FDFDFD",X"FFFCFD",X"FFFFFF",X"FEFFFF",X"FFFAFF",X"FFE7FF",X"A66689",X"3D091F",X"141C1F",X"004435",X"9FECDC",X"E3FFFF",X"FDF8FE",X"FFFBFF",X"FAFBF6",X"F6FFFC",X"F4FFFF",X"7A9793",X"3B5F5B",X"224642",X"9AB7B3",X"EDFDFA",X"F6FFFC",X"FFFAFE",X"FFFEFC",X"FFFFFD",X"FEFFFF",X"FFFEFF",X"FFFEFB",X"FFFFE1",X"FFFFC9",X"EBCC60",X"C1AF0F",X"B5AB0B",X"FFF4A4",X"FFFCF3",X"FDFBFF",X"FBFFFD",X"F6FFFF",X"FCFFFF",X"C4FFF3",X"47DBAB",X"01BF81",X"0FB881",X"A8FFF0",X"E1FFF9",X"FFFBFF",X"FAFAFA",X"FFFCFF",X"FFFBFF",X"F1F3F2",X"ECFFFB",X"B9DFD2",X"3F6055",X"000D04",X"D1C0C6",X"FFEEF6",X"FFEFF8",X"FFEAF7",X"FFE8F6",X"FFDFEF",X"FFD8E8",X"F4B4C4",X"595355",X"040000",X"070304",X"8E8A8B",X"F2F0F1",X"FFFFFF",X"FDFDFD",X"F7F9F8",X"FFFAFE",X"E9F6FF",X"658CD9",X"0D48B0",X"1651B7",X"ABD3FF",X"F2FFFF",X"FDF9EE",X"F8FFFF",X"FBF9FC",X"FFFCFF",X"FDFFFE",X"F5FFFA",X"FFFCFB",X"FFDBEC",X"B74C6A",X"AA002B",X"B03D5A",X"FFE0E5",X"F8FDF6",X"F4FEF6",X"FEFFFF",X"F5F9FA",X"F7FFFF",X"637C79",X"000606",X"010B0C",X"BBBCC0",X"FFFCFF",X"FFE9F1",X"FFE9F7",X"D29FAE",X"774455",X"FFE3F3"),
(X"EFFEFB",X"F7FFFF",X"919797",X"070105",X"070208",X"D1D5D8",X"FFFEFF",X"FDFEFF",X"FFFBFF",X"FFF2EA",X"E1DBC1",X"E7EFDA",X"FFFEFF",X"F7F6FF",X"FBFBFF",X"FFF8F9",X"FFF2FF",X"8E8A87",X"140014",X"B78EB6",X"FCEBF5",X"FFF9FD",X"FFF8FF",X"F8FFFF",X"FFFFFD",X"FFFCFE",X"FEF8FC",X"F4FDFC",X"F4FFFF",X"F4F5FF",X"E9C2F7",X"4C024F",X"E5CCE9",X"FFFAFF",X"FCF2F3",X"FEFDFF",X"FCEBFF",X"C06FB4",X"660353",X"80508A",X"E7D4EA",X"F9EAFD",X"FFFAFF",X"FFFCFF",X"FAF9FE",X"FBFCFE",X"FFFFFF",X"FDFCFF",X"FFF4FF",X"919FAA",X"040004",X"783100",X"D77826",X"FFDAB2",X"FFF8DD",X"FFFEFD",X"FFFAF0",X"FDFEF8",X"F7FEFF",X"F1F3DD",X"E0AF86",X"E48E17",X"B9711C",X"FFE3D0",X"FEFDFF",X"FEFEFF",X"FEFEFC",X"FDFFFA",X"FEFFFA",X"FEFEFC",X"FEFEFF",X"FFFDFF",X"F6FFF8",X"FFF6FF",X"EEDFE4",X"4C424D",X"100001",X"7E7854",X"F6F8ED",X"FDF4FF",X"F8FCFB",X"FFF5FF",X"D9DFEF",X"DDC5DB",X"F0F8FA",X"FBFFFD",X"FFFEFD",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FDFDFD",X"FFFFF3",X"F3DEFF",X"BD488C",X"D3006B",X"C31962",X"FFBEEA",X"FFFCEC",X"F5FFEF",X"FCEBFE",X"DE8CBD",X"C80565",X"C4005B",X"F4A7D1",X"FEF8FC",X"FFFDF8",X"F8FBF0",X"FFF0FF",X"EE7BBE",X"7E004E",X"4E153E",X"D4C8D6",X"FEFEFF",X"FBFEFF",X"FFF8FC",X"F9F8F4",X"FBFFFB",X"F5FEFB",X"FEFFFF",X"FFF6FE",X"A999A4",X"090008",X"0C1115",X"000317",X"D4DDEE",X"F4FFFF",X"F4FEFF",X"FFFCFF",X"FFF5FF",X"FAFEFF",X"9ABBC2",X"00000E",X"040100",X"5B5060",X"E9E7E8",X"FFFFEC",X"FFF6FF",X"FFFAF8",X"F7FDF1",X"FFFAFB",X"F7FDF9",X"FFFBFA",X"FFF5F9",X"837A7B",X"1B0000",X"500002",X"F99E99",X"FFF9FF",X"FFFBFF",X"FAF6F3",X"F5FBF7",X"FFFCFF",X"F2D6ED",X"21141E",X"000800",X"B1BBBA",X"FAFFFF",X"F9F9FB",X"D6D1D5",X"EEE8EC",X"FFFDFF",X"FDF7FB",X"FFFBFF",X"FFFDFE",X"F5FEFD",X"E283AB",X"C3004B",X"CC5B91",X"FCEFFF",X"FFF8FE",X"F5FFF6",X"FFFEFF",X"F9F7FA",X"C6C5CA",X"DBDCDE",X"F6F8F7",X"F8FAF9",X"FEFFFF",X"CFCED6",X"0C2C37",X"100223",X"8295A4",X"F1FAFF",X"FFF3F9",X"F9FDFE",X"EDFEFF",X"CAE5EE",X"C5D8DF",X"FCFFFF",X"EFFFFF",X"F5FFF6",X"FFF7F6",X"DFFFFF",X"6AD5FF",X"00567A",X"000606",X"C1BEB9",X"FFFCF4",X"FFF7F3",X"FFFEFF",X"F7FCFF",X"F8FEFE",X"FEFFFA",X"FEFDF9",X"F7FFFF",X"FCFFF4",X"FEF5D4",X"B6AD8C",X"6B6E63",X"F9FEFF",X"FFFAFE",X"F8FBF0",X"F9FFF4",X"FBC5DC",X"CF3275",X"B40349",X"C56298",X"FEECFF",X"F7FEF6",X"FFFFFF",X"FDF6FD",X"FEFFFF",X"FAFCFB",X"FFFDFD",X"FFFDFE",X"FFF0FC",X"DF99BE",X"2D0304",X"110000",X"24413C",X"C2E2DF",X"FCF2FA",X"FFF5FA",X"F9FFFD",X"F7FFFD",X"FCFCFF",X"E5FDFF",X"78B5B0",X"08AB8E",X"38B1AA",X"079B8B",X"84DDD9",X"D8FFFF",X"F2FFFF",X"F1FFFB",X"F3FFF5",X"FBFEF7",X"FFFAFE",X"FAF7FE",X"FEFFFF",X"F8FBF2",X"F3DF9A",X"BBA600",X"D2B245",X"FFF4D6",X"FFFFFD",X"FBF9FF",X"FFFFF1",X"FAF7FE",X"FBFFF9",X"F3F7F8",X"86C0B2",X"32B394",X"37AD7D",X"D8F3FC",X"FFFDF2",X"F7FFFE",X"FAF8F9",X"F9FFFF",X"FFEEF9",X"EFFFFF",X"91FFE6",X"00B280",X"44A287",X"C9DAD2",X"FEFDFB",X"FFFCFD",X"FFF9FE",X"FFF8FF",X"FEF9FF",X"FEF9FD",X"FFF8FC",X"FFF8FB",X"E8DCE6",X"443E42",X"1A1914",X"010700",X"9DA097",X"FFF8F6",X"FCF8F9",X"F2FFFF",X"FFFCFF",X"FAFBEB",X"91AFE1",X"002EAC",X"225AB9",X"CFDEF1",X"FFFEF8",X"F7FFFF",X"FFFCFF",X"F7FFF4",X"FBFFF6",X"FFF8FF",X"FFFCFF",X"FAFFFB",X"FBEDED",X"BE8DA2",X"890007",X"C27484",X"F6E4F0",X"FFFFFD",X"FFFEFF",X"F6F8FF",X"FCFEFF",X"FFFCFF",X"BD889A",X"560000",X"2E0005",X"E0CFDF",X"FFFAF8",X"FFFAFB",X"F4FFF6",X"FFF5FF",X"D3C5C5",X"FEF6F4"),
(X"F5FFFF",X"F2FEFC",X"B1B7B7",X"090307",X"030004",X"DDE1E4",X"FCFBFF",X"FCFDFF",X"FAEEF2",X"FFF8F0",X"FFFBE1",X"FCFFEF",X"FDFBFF",X"FBFAFF",X"F7F7FF",X"FFF8F9",X"C6AFBF",X"050100",X"856D85",X"FFDCFF",X"FFF5FF",X"FFF3F7",X"FFF9FF",X"F8FFFF",X"FCFCFA",X"FFFCFE",X"FFFDFF",X"EFF8F7",X"EDFCFF",X"FCFDFF",X"FCD5FF",X"540A57",X"DCC3E0",X"FDF1FB",X"FFFCFD",X"FBFAFF",X"B7A6C6",X"550449",X"832070",X"F4C4FE",X"FFEFFF",X"FFF5FF",X"FFFAFF",X"FFFCFF",X"FEFDFF",X"FEFFFF",X"FEFEFF",X"FCFBFF",X"FFF6FF",X"EDFBFF",X"867F86",X"9A5313",X"DD7E2C",X"D39E76",X"FFFFE4",X"F8F4F3",X"FFFEF4",X"F9FAF4",X"F5FCFF",X"F9FBE5",X"D2A178",X"D07A03",X"F1A954",X"FFDECB",X"FEFDFF",X"FEFEFF",X"FEFEFC",X"FDFFFA",X"FEFFFA",X"FEFEFC",X"FEFEFF",X"FFFDFF",X"F9FFFB",X"FFF2FF",X"F6E7EC",X"625863",X"0D0000",X"BDB793",X"FFFFF6",X"FBF2FF",X"F8FCFB",X"FFF3FF",X"F7FDFF",X"FFF2FF",X"F7FFFF",X"F8FEFA",X"FFFBFA",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FDFDFD",X"FFFBEF",X"FAE5FF",X"E36EB2",X"C7005F",X"D42A73",X"FFBEEA",X"FFFFEF",X"EEFDE8",X"FFF6FF",X"FFB8E9",X"CB0868",X"CE0565",X"BC6F99",X"FAF4F8",X"FFF6F1",X"FEFFF6",X"E8CDDE",X"932063",X"951665",X"E1A8D1",X"FFFAFF",X"F8F8FF",X"F4F7FE",X"FFFAFE",X"FDFCF8",X"FAFFFA",X"F9FFFF",X"F6F7F9",X"FEF4FC",X"FFF6FF",X"9B919A",X"04090D",X"000013",X"5D6677",X"E3F1FA",X"F4FEFF",X"FFFBFF",X"FFF5FF",X"FBFFFF",X"B6D7DE",X"050716",X"040100",X"736878",X"F5F3F4",X"FFFCE9",X"FFF0F9",X"FFFAF8",X"FCFFF6",X"FEF5F6",X"FBFFFD",X"FFFBFA",X"FEF2F6",X"E6DDDE",X"4D2629",X"59070B",X"A34843",X"EFE7F4",X"FFF9FD",X"FFFEFB",X"F9FFFB",X"FFFDFF",X"C8ACC3",X"0A0007",X"7F9588",X"F4FEFD",X"FBFFFF",X"FFFFFF",X"FFFAFE",X"FFF9FD",X"FFF9FD",X"FFF9FD",X"FFFAFE",X"FFFBFC",X"F6FFFE",X"E687AF",X"C90051",X"D16096",X"FEF1FF",X"FFF8FE",X"F3FFF4",X"FDFBFC",X"FFFEFF",X"F4F3F8",X"FCFDFF",X"FEFFFF",X"FAFCFB",X"FEFFFF",X"E3E2EA",X"365661",X"060019",X"738695",X"F8FFFF",X"FFF1F7",X"FCFFFF",X"E8F9FF",X"E6FFFF",X"ECFFFF",X"F2F5FC",X"F1FFFF",X"F9FFFA",X"FFF6F5",X"C1E4FF",X"1F8AB6",X"1082A6",X"B3B9B9",X"FFFFFA",X"FFFCF4",X"FDF2EE",X"FEFCFF",X"F6FBFF",X"FBFFFF",X"FEFFFA",X"FEFDF9",X"F7FFFF",X"F0F6E8",X"FFFFDF",X"CCC3A2",X"717469",X"F3F8FC",X"FFFDFF",X"FAFDF2",X"F8FFF3",X"FFD5EC",X"D93C7F",X"B30248",X"D976AC",X"FFF5FF",X"F9FFF8",X"FDFDFF",X"FFF9FF",X"FDFEFF",X"FDFFFE",X"FCF6F6",X"FDFBFC",X"FFF8FF",X"FFBEE3",X"270000",X"0F0000",X"203D38",X"CBEBE8",X"FFFBFF",X"FFF7FC",X"F8FFFC",X"F1FEF7",X"F9F9FF",X"E9FFFF",X"79B6B1",X"0BAE91",X"2DA69F",X"1EB2A2",X"27807C",X"9ECED0",X"F4FFFF",X"E6FCF0",X"F4FFF6",X"FCFFF8",X"FFFDFF",X"FFFDFF",X"F8FAF9",X"FEFFF8",X"F1DD98",X"B49F00",X"D4B447",X"FFF5D7",X"FEFEFC",X"FCFAFF",X"FFFFF1",X"FFFCFF",X"F6FBF4",X"FCFFFF",X"75AFA1",X"005D3E",X"108656",X"DCF7FF",X"FFFBF0",X"F6FFFD",X"FFFEFF",X"EFF8F5",X"FFF6FF",X"E0F6F4",X"37A88C",X"00AA78",X"86E4C9",X"EFFFF8",X"FDFCFA",X"FFFBFC",X"FFF9FE",X"FFF9FF",X"FFFAFF",X"FEF9FD",X"FFF7FB",X"FFF6F9",X"FFFAFF",X"C8C2C6",X"010000",X"1F2519",X"020500",X"EBE3E1",X"FAF6F7",X"F4FFFF",X"FFFCFF",X"FFFFF1",X"98B6E8",X"003AB8",X"3169C8",X"D6E5F8",X"FFFEF8",X"F9FFFF",X"FFFDFF",X"F7FFF4",X"FBFFF6",X"FFF9FF",X"FFFCFF",X"FBFFFC",X"FFF4F4",X"CC9BB0",X"870005",X"CF8191",X"FEECF8",X"FDFDFB",X"FFFEFF",X"F8FAFF",X"FCFEFF",X"FFFCFF",X"DCA7B9",X"6E110A",X"58172F",X"D9C8D8",X"FFFAF8",X"FFFCFD",X"F6FFF8",X"FFF4FF",X"FFFBFB",X"FFFDFB"),
(X"F7FBFC",X"FFF7FE",X"B8B8BA",X"000F07",X"000004",X"F3D9E6",X"FDFBFF",X"F6FAFD",X"F1FFFF",X"FEFBFF",X"FFFCFF",X"F9F9FB",X"FCF8F9",X"FBFFFF",X"F5FEFF",X"F7ECFC",X"5D287A",X"170028",X"D7B9DD",X"FFFBFF",X"F6FFF9",X"FBFFFF",X"FFFDFF",X"FAFBF3",X"F6FFFF",X"FAFDFF",X"FFFAFE",X"FFFAFA",X"FFF9F6",X"FFF5F4",X"FDF4F9",X"BDBAC5",X"FFEBFF",X"F5FFFF",X"F6FFFC",X"EBDEE7",X"633E5D",X"4C0E3F",X"D6A1CD",X"FFF9FF",X"FFFEFF",X"FEFEFC",X"FBFDF8",X"FBFFF9",X"FCFFFA",X"FEFFFB",X"FEFEFC",X"FEFEFE",X"FCF6F8",X"FCFFF8",X"F1E4DB",X"C8824F",X"F7861C",X"DF8515",X"FFE0A1",X"FFF9FF",X"F2F8FF",X"F6F0F4",X"FFFEFF",X"FFFEFA",X"B7A6B8",X"150000",X"A1856D",X"FFF0E9",X"FFF9FF",X"FFFAFF",X"FFFBFF",X"FFFCFF",X"FFFDFE",X"FFFDFE",X"FEFEFE",X"FEFEFE",X"FBFFF8",X"FFFFF4",X"EAF6F4",X"64686B",X"7F6E28",X"D5C868",X"FFFFEC",X"F8FFF7",X"FAFFF1",X"FFF2F9",X"FAF8FF",X"FFFCFF",X"F8FFF8",X"FFFEFF",X"FFFDFF",X"FCFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FDFDFD",X"F5FFF8",X"FFE8FF",X"E771A3",X"C21161",X"C6488F",X"FFD7FF",X"FFF3FF",X"FFF7FF",X"FDF9FF",X"FFDFF2",X"D26491",X"8D1147",X"AB7899",X"FFF7FF",X"FFF3FF",X"F5F9FA",X"957584",X"530F26",X"8E5F69",X"EEF0E5",X"F3FDF4",X"F6FBF7",X"FDFFFA",X"FFFEF6",X"FFFDFF",X"F9F2F9",X"FFF6FF",X"FFF9FF",X"F5FDFF",X"FFFCFF",X"FFECF8",X"807B81",X"080007",X"000013",X"AFBAD6",X"FCFBFF",X"FFFEFB",X"F8FFF1",X"F4FCFE",X"DFD9F3",X"263560",X"000300",X"857F8B",X"F9FBFF",X"F9FFFD",X"FDFAFF",X"FDFCFA",X"F7FFFF",X"FEFEFE",X"FCFBF9",X"FAFFFE",X"F3FFFF",X"FAFEFD",X"D9B1B9",X"710817",X"A00018",X"F68D91",X"FFEFF7",X"FEFCFF",X"FFF4F0",X"FFE3DA",X"9A394D",X"621E35",X"E4EAEA",X"F9FFFF",X"F0F4F5",X"F8F8FA",X"FFFDFF",X"FCF6FA",X"FEF8FC",X"FFFDFF",X"FBF9FC",X"FAF9FF",X"F9FCFF",X"EB86B0",X"CD0253",X"D76098",X"FFF2FF",X"FFF9FF",X"F5FFF9",X"F9F7F8",X"FCFCFE",X"FFFEFF",X"FDFEFF",X"F9FBF8",X"FCFCFA",X"FBF9FE",X"F1EEF7",X"9B5480",X"2A0004",X"8A837D",X"F5F9FA",X"EEFDF8",X"F4FFF1",X"FFF5F0",X"FFF7FF",X"FEFDF8",X"FFFAFF",X"FEFFFF",X"FFFFF1",X"DEF7FC",X"5DD4FF",X"0695D7",X"70A2C3",X"EDFFFF",X"F7FFFF",X"FAFBFD",X"FEFCFF",X"FFFDFF",X"FCFAFF",X"FFFAFF",X"FFF5FE",X"FFFCFA",X"FBFCFF",X"FFFFFD",X"FFFEEF",X"F1E8D9",X"C5C5C5",X"FFFEFF",X"FFF8FA",X"FFF8FF",X"F7FFFF",X"F2F5FF",X"876371",X"4A151D",X"AB8E93",X"FCF5FC",X"FFFAFE",X"FCFFFA",X"FFFEFF",X"F9FEFF",X"FBFFFF",X"FFFEFF",X"F8FFFF",X"FFFCFD",X"F5C5D5",X"57000C",X"220509",X"2D443E",X"D3E9E6",X"F8FFFF",X"F6FAF9",X"FFFDFE",X"FFF9FF",X"FFFCFF",X"DEFEF9",X"65BEAA",X"00B488",X"21BB9F",X"0FAC8F",X"1EA489",X"009670",X"7CE7D5",X"E2FFFF",X"FFF7FF",X"FEFEFF",X"F1FDFD",X"FCF5FC",X"FFFCFB",X"F3FFEF",X"F5E6AD",X"B69708",X"DABB6B",X"FFFFE8",X"F8FFF7",X"FDF9FF",X"FFFEFA",X"FFFFF6",X"FAFEFF",X"FFFBF9",X"A5A38E",X"000F00",X"565D33",X"F7E3EF",X"FFFBF8",X"F9FEFF",X"FFFDFF",X"EFFBF7",X"FEFFFF",X"AACAC5",X"17A17D",X"38C09C",X"C6FAED",X"F8FCFB",X"F5FDFF",X"F7FCFF",X"F9FCFF",X"F9FEFF",X"F6FFFF",X"F5FFFF",X"F7FCFF",X"FAF9FE",X"FAFCF7",X"F5FAFF",X"947A95",X"1B0012",X"040007",X"8B868A",X"FFF9FF",X"FBF5FF",X"FDF8FF",X"FFFEF7",X"9FB6DF",X"053BA8",X"3A6FCD",X"D2E4FC",X"FFFFFA",X"F8FBFF",X"FFFBFF",X"FAFDFF",X"F9FFFF",X"FCFDF8",X"FEFFF7",X"FCFDF7",X"FFF6FC",X"E2A9BC",X"7D0002",X"D894A1",X"FFF5FF",X"FAF9FE",X"FFFCFC",X"FFFCFF",X"FCFFFF",X"FCFFF4",X"EAC1BD",X"740000",X"9D2D51",X"F9D7E5",X"FFF8EF",X"FEF9FF",X"F5FFFF",X"F8FFFF",X"FFF2F9",X"FDF7FB"),
(X"FCFFFF",X"FFFAFF",X"D3D3D5",X"000A02",X"040308",X"E1C7D4",X"FFFEFF",X"FAFEFF",X"EDFFFF",X"F9F6FF",X"FFFDFF",X"FBFBFD",X"FFFEFF",X"F6FCFC",X"F5FEFF",X"C9BECE",X"3A0557",X"471E58",X"D3B5D9",X"FFFBFF",X"F4FFF7",X"F1F7F7",X"FFFDFF",X"FBFCF4",X"F3FDFF",X"FCFFFF",X"FFFAFE",X"FFF9F9",X"FFFBF8",X"FFF6F5",X"FFF8FD",X"FFFDFF",X"FFECFF",X"EFFDFF",X"F7FFFD",X"C0B3BC",X"160010",X"2E0021",X"FFCAF6",X"FFF7FF",X"FBF9FA",X"FCFCFA",X"FEFFFB",X"FCFFFA",X"FBFFF9",X"FCFEF9",X"FEFEFC",X"FFFFFF",X"FFFAFC",X"F2F8EE",X"FFFBF2",X"F5AF7C",X"EF7E14",X"E28818",X"D0AE6F",X"FFFBFF",X"F9FFFF",X"FFFDFF",X"F2F0F3",X"FFFEFA",X"CFBED0",X"110000",X"866A52",X"FFF2EB",X"FFF9FF",X"FFFAFF",X"FFFBFF",X"FFFCFF",X"FFFDFE",X"FFFDFE",X"FEFEFE",X"FEFEFE",X"F8FFF5",X"F9FBEE",X"F7FFFF",X"6C7073",X"85742E",X"F0E383",X"F8FAE4",X"EFF6EE",X"F9FFF0",X"FFFAFF",X"FBF9FF",X"F9F3F7",X"FBFFFB",X"FFFEFF",X"FCF7FD",X"FCFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FDFDFD",X"F6FFF9",X"FFEDFF",X"F07AAC",X"AE004D",X"C5478E",X"FFDBFF",X"FFF0FF",X"FFF6FF",X"FFFCFF",X"FFE6F9",X"D0628F",X"74002E",X"D29FC0",X"FAEDFF",X"FFF8FF",X"CDD1D2",X"190008",X"2D0000",X"A67781",X"FBFDF2",X"F8FFF9",X"FCFFFD",X"F7F9F4",X"FFF9F1",X"FFFAFE",X"FFFCFF",X"FFF4FE",X"FFFBFF",X"F9FFFF",X"FAF3FB",X"FFF7FF",X"C0BBC1",X"090008",X"000518",X"77829E",X"F4F3FF",X"FDF8F5",X"FBFFF4",X"F9FFFF",X"F1EBFF",X"51608B",X"000400",X"938D99",X"F9FBFF",X"F9FFFD",X"FFFDFF",X"FDFCFA",X"F2FCFE",X"FFFFFF",X"FEFDFB",X"F8FEFC",X"F4FFFF",X"F8FCFB",X"FFEDF5",X"D16877",X"9E0016",X"A73E42",X"F8E1E9",X"FFFDFF",X"FFF5F1",X"D7ABA2",X"67061A",X"FEBAD1",X"F5FBFB",X"F3FCFB",X"FCFFFF",X"FDFDFF",X"FAF5F9",X"FCF6FA",X"FFFAFE",X"FFFBFF",X"FDFBFE",X"FCFBFF",X"F9FCFF",X"E984AE",X"C9004F",X"D25B93",X"FDEFFF",X"FFF9FF",X"F7FFFB",X"FEFCFD",X"FAFAFC",X"FCFBFF",X"F8F9FB",X"F9FBF8",X"FFFFFD",X"FFFEFF",X"F8F5FE",X"B06995",X"480F22",X"938C86",X"FAFEFF",X"F5FFFF",X"EAFDE7",X"FFFBF6",X"FFF8FF",X"FDFCF7",X"FFF9FF",X"F2F3F7",X"FFFFF1",X"D4EDF2",X"188FC7",X"0F9EE0",X"92C4E5",X"ECFFFF",X"EEF9FF",X"FBFCFE",X"FFFDFF",X"F9F7FF",X"FCFAFF",X"FFFBFF",X"FFF9FF",X"FFF9F7",X"F9FAFE",X"FFFFFD",X"FFF6E7",X"FFFCED",X"FFFFFF",X"FFFEFF",X"FCF0F2",X"FEF0FF",X"F3FBFF",X"F0F3FF",X"724E5C",X"240000",X"9E8186",X"FFFCFF",X"FEF9FD",X"F9FEF7",X"FFFEFF",X"FBFFFF",X"F9FDFF",X"FEFDFF",X"F1FBFA",X"FFFCFD",X"FFD1E1",X"520007",X"1A0001",X"3B524C",X"DCF2EF",X"F8FFFF",X"FBFFFE",X"FFFEFF",X"FFF7FD",X"FFFCFF",X"E9FFFF",X"5EB7A3",X"009F73",X"3BD5B9",X"2ECBAE",X"088E73",X"13A983",X"26917F",X"C3E1E1",X"FFEEF6",X"FFFFFF",X"F7FFFF",X"FFFBFF",X"FFF9F8",X"F8FFF4",X"FEEFB6",X"B69708",X"E1C272",X"FFFFEA",X"F6FDF5",X"FEFAFF",X"FCFBF7",X"FEFEF4",X"FCFFFF",X"FAF2F0",X"BFBDA8",X"47561F",X"80875D",X"FCE8F4",X"FFFBF8",X"FAFFFF",X"FDF7F9",X"F5FFFD",X"F7F9F8",X"54746F",X"17A17D",X"4ED6B2",X"D4FFFB",X"F9FDFC",X"F6FEFF",X"F8FDFF",X"FAFDFF",X"F9FEFF",X"F6FFFF",X"F5FFFF",X"F8FDFF",X"FBFAFF",X"FAFCF7",X"FBFFFF",X"D7BDD8",X"350C2C",X"09010C",X"3E393D",X"E9D8E2",X"FFFCFF",X"FEF9FF",X"FFFFF8",X"A4BBE4",X"053BA8",X"3A6FCD",X"D1E3FB",X"FFFFFA",X"FBFEFF",X"FFFBFF",X"F9FCFF",X"F9FFFF",X"FDFEF9",X"FCFDF5",X"F9FAF4",X"FFF7FD",X"EBB2C5",X"7C0001",X"E4A0AD",X"FFF8FF",X"F8F7FC",X"FFFDFD",X"FFFDFF",X"FAFEFD",X"FDFFF5",X"EBC2BE",X"820A0B",X"A9395D",X"FDDBE9",X"FFFBF2",X"FFFDFF",X"F5FFFF",X"F2F9FF",X"FFFAFF",X"FFFBFF"),
(X"FFF5FB",X"FCFCFE",X"C3E1D9",X"001602",X"000306",X"FCDCEB",X"FAFEFF",X"FFECFB",X"FFEDFF",X"FFE0FF",X"FFD8FF",X"FFEEFF",X"FFFAF9",X"F9F9EF",X"FFF7FF",X"AF7DAE",X"74007F",X"79067F",X"EBA9E7",X"FFFAFA",X"FCFFFF",X"FCF6FF",X"FDFEFF",X"F5FFEF",X"FFFCFA",X"FFFCF9",X"FBFFFD",X"F9FFFA",X"F5FBF1",X"FFFFF8",X"FFFFFD",X"F7F5FA",X"FFF6FF",X"FFF9FF",X"F8F4F5",X"4F5B5B",X"00120E",X"000D0B",X"D1DFE0",X"FFFFFB",X"FAF9F4",X"FFFFF8",X"FFFFF8",X"FFFFFA",X"FFFCF9",X"FFFBFB",X"FFFAFE",X"FFF8FF",X"F7FFFF",X"FFFDFF",X"FFFCF0",X"FCD39F",X"E87300",X"F17400",X"E0A374",X"FFFCEC",X"EEF9FF",X"FAEFF7",X"FEFFFB",X"FDF4F7",X"C1C8FE",X"000B66",X"717D97",X"F2F7F3",X"F7FFF2",X"F7FFF3",X"F8FFF7",X"FAFFFA",X"FBFFFC",X"FDFFFE",X"FEFEFE",X"FFFDFE",X"F5FFFF",X"F9FFF1",X"F6FFFC",X"7F7F87",X"53460F",X"E1D99B",X"F8F3FA",X"FFFAFF",X"FEF5F6",X"FFF2FF",X"FFDEFF",X"FFFDFF",X"FEFFF8",X"FFFEFF",X"FFFCFF",X"FEFFFD",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FDFDFD",X"FDFCFF",X"FFF9FF",X"C697A9",X"531522",X"855D7F",X"FCEAF6",X"FFF5EF",X"FFFBF0",X"FAF6F3",X"CDD6D1",X"1B040C",X"1B0002",X"E7DAE3",X"FFFBFF",X"FFF8FF",X"ADC2DF",X"000C2E",X"000427",X"96A2BA",X"FCFFFF",X"FFF4F4",X"FFF9F5",X"FAFFF9",X"F9FFFB",X"F6FFFB",X"FCFFFD",X"FFF9FA",X"FFFDFD",X"F4FFF9",X"FFFFFB",X"FFFEFA",X"C7D5C8",X"363835",X"07000E",X"0A0022",X"D1DDED",X"F5FFFD",X"FBF9ED",X"FEF3F7",X"F4F1FF",X"4D68AF",X"000209",X"9F9697",X"FEFCFF",X"F1FAFF",X"F8FDFF",X"FCFEF9",X"FBFFFF",X"F1FFFB",X"FFF9FF",X"FFF9FD",X"FCFFFF",X"FFFCFF",X"FEEFF4",X"FFD9DF",X"A53647",X"A10000",X"FF779A",X"FFE0F7",X"FFD4D4",X"8E060A",X"B67476",X"ECF2F0",X"FFF2FD",X"F9FDFE",X"FEFFFF",X"FFFEFF",X"FFFAFE",X"FFFDFF",X"FFFCFF",X"F9F9FB",X"FFFFFF",X"FAFDFF",X"FDFAFF",X"E385AA",X"BF0048",X"D05A8E",X"FBEFFD",X"FFFCFF",X"F9FFFF",X"FCFCFC",X"FFFFFF",X"FFFEFF",X"FFFFFF",X"FFFFFD",X"FFFEFC",X"FFFDFF",X"F7EFFA",X"CD5C92",X"8C154B",X"AE8299",X"FEFFFF",X"F1F8FF",X"DEFFFF",X"D3FFFF",X"E1FCFF",X"EBFAFF",X"FFF5F8",X"FFFDF4",X"FEFFFD",X"C5E6FF",X"0088D9",X"00A4E4",X"B0E0F7",X"FFFFFF",X"FFFEFB",X"FFFFF6",X"F9FBF0",X"F6FDF5",X"F8FFFB",X"F8FFF8",X"FBFFF6",X"FFFBF8",X"FFFEFF",X"F9FAFF",X"FFF9F9",X"FFFDFD",X"F8FBFF",X"FEFFFF",X"FFFBF8",X"FFFBFA",X"F4F8F9",X"F5FFED",X"AFC16D",X"4A5300",X"959639",X"FCFDC3",X"FFFFD3",X"F8FFD1",X"FFFCE3",X"FEEEEE",X"FFECFF",X"FFDBFF",X"FFDEFF",X"FFD1FF",X"FFA6E4",X"7C082D",X"1D0007",X"5A595E",X"FDF4F9",X"FAFFFB",X"F8FFFD",X"FFFBFF",X"FFFBFF",X"FFFBFE",X"E8F8F5",X"89B4AB",X"317B6C",X"8ECDC4",X"D4FCFB",X"63A297",X"119973",X"0EAA92",X"209F8A",X"A7F9EB",X"DDFFFC",X"FEFFFF",X"FFF9FF",X"FFF5F3",X"FFFFF3",X"F8EDB5",X"B69102",X"DCC174",X"F6FFF2",X"F3FFF5",X"FFFBFF",X"FCFCFE",X"FEFFF5",X"FFFBFF",X"FCF8EF",X"DCCB97",X"C2A82F",X"C6A764",X"FFF8F5",X"FCFAFB",X"FFFBFF",X"F9FDFC",X"F4FFFF",X"C1C5C4",X"000104",X"30A185",X"94DECF",X"E2F4F4",X"F8FFFE",X"FFFFFA",X"FFFDFA",X"FFFCFC",X"FEFDFB",X"FCFEFB",X"FAFFFB",X"FEFFFA",X"FFFEF9",X"FFFEFA",X"EEFFFF",X"F6E5FF",X"CA5FAF",X"890F64",X"2D0025",X"D6C5D8",X"FFFAFF",X"FBF9FF",X"FFFDFF",X"B6C1D7",X"0A3480",X"3563B9",X"CADFFC",X"FFFFFA",X"FFFBFF",X"FFFBFF",X"FAFAFF",X"FBFFFF",X"FBFFF7",X"FCFFF6",X"FAF7FE",X"FFF6FF",X"E9B9B5",X"5E0700",X"DAADB2",X"FFFAFF",X"FAF9FE",X"FFFCFD",X"FFFDFF",X"FAFCF7",X"FBFFF6",X"F7C8DC",X"8C000C",X"D34462",X"FFE3F3",X"FFF1F8",X"FFE4F6",X"FFE7F1",X"FFE1F1",X"F8EBF5",X"FFFBFF"),
(X"FFF5FB",X"FFFFFF",X"D4F2EA",X"11523E",X"000104",X"C5A5B4",X"D1D5D8",X"C5A5B4",X"A37E9D",X"9D6596",X"875B8E",X"EEDCF6",X"FFF8F7",X"FDFDF3",X"FFF3FF",X"A16FA0",X"770382",X"7E0B84",X"F4B2F0",X"FCF6F6",X"F9FDFC",X"FFFCFF",X"F6F7F9",X"F5FFEF",X"FFFCFA",X"FFFDFA",X"FBFFFD",X"F9FFFA",X"FAFFF6",X"FEFFF7",X"FFFEFC",X"FFFEFF",X"FFF3FF",X"FFFAFF",X"F4F0F1",X"3B4747",X"315B57",X"1E4846",X"D7E5E6",X"FFFFFB",X"FDFCF7",X"FFFFF8",X"FFFFF7",X"FCFBF6",X"FFFBF8",X"FFFDFD",X"FFFBFF",X"FFF7FE",X"F4FEFF",X"FFFBFD",X"FFFFF3",X"FFDBA7",X"F6810D",X"EC6F00",X"E9AC7D",X"FFFAEA",X"F5FFFF",X"FFF5FD",X"FBFDF8",X"FFFCFF",X"BCC3F9",X"0E338E",X"6E7A94",X"F6FBF7",X"F7FFF2",X"F7FFF3",X"F8FFF7",X"FAFFFA",X"FBFFFC",X"FDFFFE",X"FEFEFE",X"FFFDFE",X"F5FFFF",X"FAFFF2",X"F8FFFE",X"818189",X"130600",X"91894B",X"D9D4DB",X"C3B4BB",X"A39A9B",X"917792",X"8F5F85",X"E0DADE",X"F6F9F0",X"FDFBFE",X"FFFDFF",X"F4F6F3",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FDFDFD",X"FCFBFF",X"FFFAFF",X"B28395",X"2A0000",X"684062",X"FFF0FC",X"FFFCF6",X"FFF9EE",X"FBF7F4",X"636C67",X"110002",X"D4ABBB",X"FFFAFF",X"F9F1FF",X"FEF3FF",X"8CA1BE",X"0E4466",X"2B4568",X"C4D0E8",X"FCFFFF",X"FFF4F4",X"FFFCF8",X"FBFFFA",X"EDF7EF",X"F8FFFD",X"F7FCF8",X"FFF5F6",X"FFFDFD",X"F0FBF5",X"FBFCF7",X"FFFEFA",X"F5FFF6",X"494B48",X"0C0013",X"03001B",X"CBD7E7",X"F3FFFB",X"FDFBEF",X"FFFBFF",X"F7F4FF",X"4D68AF",X"000209",X"A09798",X"FFFDFF",X"F4FDFF",X"F7FCFF",X"FCFEF9",X"FBFFFF",X"F5FFFF",X"FFF8FE",X"FFFAFE",X"FCFFFF",X"FCF7FD",X"FFF7FC",X"FFECF2",X"F38495",X"A90000",X"94082B",X"F2BED5",X"CA8484",X"8D0509",X"FFD0D2",X"F7FDFB",X"FFF2FD",X"FAFEFF",X"F9FAFC",X"FDFBFE",X"FFFDFF",X"FFFDFF",X"FFFDFF",X"FFFFFF",X"FEFEFF",X"FBFEFF",X"FDFAFF",X"E385AA",X"C00049",X"D25C90",X"FDF1FF",X"FFFCFF",X"F8FFFE",X"FCFCFC",X"FFFFFF",X"FAF9FE",X"FFFFFF",X"FFFFFD",X"FBFAF8",X"FFFDFF",X"F2EAF5",X"D6659B",X"6C002B",X"8E6279",X"D5D6DA",X"BFC6D0",X"A3CDD9",X"8ABECB",X"7D98A9",X"C2D1D6",X"FFFAFD",X"FEFAF1",X"F3F5F2",X"B2D3FE",X"0697E8",X"00A0E0",X"9FCFE6",X"FAFAFC",X"FFFCF9",X"FFFDF4",X"FCFEF3",X"FBFFFA",X"F8FFFB",X"F2FEF2",X"FAFFF5",X"FFFDFA",X"FFFEFF",X"FEFFFF",X"FFFDFD",X"FFFDFD",X"F9FCFF",X"FAFBFF",X"FFFEFB",X"FFFBFA",X"FCFFFF",X"E5F7DD",X"D4E692",X"D2DB68",X"BFC063",X"BDBE84",X"DCDFB0",X"C6CE9F",X"685E45",X"160606",X"54344B",X"6C385E",X"724066",X"74305F",X"9B2967",X"982449",X"24030E",X"58575C",X"FDF4F9",X"F9FEFA",X"F6FFFB",X"FEF9FD",X"FFFCFF",X"FEF5F8",X"F4FFFF",X"6A958C",X"001A0B",X"73B2A9",X"E3FFFF",X"B8F7EC",X"33BB95",X"09A58D",X"179681",X"37897B",X"C1E4E0",X"F8F9FE",X"FFF6FD",X"FFFCFA",X"F9F7EA",X"F8EDB5",X"BD9809",X"DEC376",X"F6FFF2",X"F5FFF7",X"FFFBFF",X"FDFDFF",X"FFFFF6",X"FEF9FF",X"FFFFF6",X"DBCA96",X"BDA32A",X"D0B16E",X"FDEFEC",X"FFFEFF",X"FFFCFF",X"F6FAF9",X"EFFFFA",X"C2C6C5",X"000104",X"0D7E62",X"8DD7C8",X"F0FFFF",X"F7FFFD",X"FFFFFA",X"FFFEFB",X"FFFCFC",X"FEFDFB",X"FCFEFB",X"FBFFFC",X"FFFFFB",X"FFFFFA",X"FEF9F5",X"EDFFFF",X"F9E8FF",X"DB70C0",X"A42A7F",X"3C0034",X"DCCBDE",X"FFFAFF",X"F9F7FF",X"FFFBFD",X"BEC9DF",X"002975",X"214FA5",X"C4D9F6",X"FDFEF8",X"FCF8FF",X"FFF9FD",X"F9F9FF",X"FBFFFF",X"FBFFF7",X"FEFFF8",X"FDFAFF",X"FFF6FF",X"E7B7B3",X"540000",X"D8ABB0",X"FFF9FF",X"FCFBFF",X"FFFCFD",X"FFFCFE",X"F9FBF6",X"FBFFF6",X"F3C4D8",X"950415",X"C53654",X"ECB7C7",X"DCC7CE",X"B2899B",X"AB7D87",X"804B5B",X"B4A7B1",X"F7F0F8"),
(X"FFFBFF",X"FFFDFF",X"BFF4E4",X"00B67A",X"007147",X"000104",X"010004",X"361C29",X"582045",X"49043B",X"441448",X"F5E3FB",X"FFFEFA",X"FFFDF1",X"FFE8FA",X"B06CA7",X"8C057E",X"860085",X"EBA8EB",X"F8FFF3",X"F3F6ED",X"FFF3FF",X"FFF8FF",X"F8FFFF",X"F3FDF4",X"FFFFFD",X"FFFBFF",X"F8F6FB",X"F9FFFF",X"F8FFFF",X"F9F7FF",X"FDF0FF",X"F9FFFF",X"FDF6FD",X"E2F9F3",X"48BE9C",X"26E9AF",X"22CF9A",X"BBFFEB",X"FBFDF2",X"F6FEFF",X"F5FDFF",X"F6FBFE",X"F8FCFF",X"FBFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"F9FFFF",X"FEF5FF",X"F7FFFF",X"FAE7BF",X"FF9126",X"EA690B",X"CC9181",X"FDF8E2",X"F4F8F7",X"FFFAFE",X"F2FFFB",X"FDF6EC",X"B5C7EB",X"0344BA",X"6C8AB0",X"EBFBFB",X"FAFFFF",X"FBFEFF",X"FBFEFF",X"FDFDFF",X"FDFDFF",X"FDFEFF",X"FDFFFC",X"FDFFF9",X"FCFFFF",X"FEF9F3",X"FFFFF4",X"9B8792",X"180009",X"150008",X"070007",X"23051F",X"0B0012",X"290136",X"5E044A",X"FDECFE",X"FFFFFB",X"F5F9FC",X"FEFFFF",X"FFFFFA",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FDFDFD",X"FCF7FB",X"FFFFFA",X"A9A781",X"0B0A00",X"66632E",X"EDF2BC",X"FEFDCF",X"E2E2A2",X"655442",X"000400",X"A0A8B3",X"E1E0E5",X"FAFFF0",X"FAFFF5",X"E7F3FF",X"6896C7",X"1175D3",X"1869C4",X"A1CFFF",X"F1FBFF",X"FFFBF4",X"FFFEFF",X"FBFCFF",X"FFFBFF",X"FFF8FB",X"FFFCFD",X"FCFEFD",X"FBFFFF",X"FFFFFF",X"FEFFFF",X"FDF7F7",X"FFEAF2",X"774F50",X"0E0000",X"030002",X"D5D2D9",X"FFFDFF",X"FAFBFF",X"FBFFFF",X"EAEFF3",X"4A6DBF",X"00011E",X"9F908D",X"FFFCFA",X"FCFFFF",X"FEFFFF",X"FFFEF9",X"FFFAFE",X"F2FFFF",X"FFFAFE",X"FFF3F9",X"FFF7FF",X"FFFDFF",X"EFF9FA",X"F8FFFB",X"EAE1DA",X"A81424",X"A8001B",X"D22E46",X"A00314",X"D8898C",X"FBF7F6",X"FEEFF6",X"F2FFF4",X"FEFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FDFBFE",X"FFFFFF",X"FEFFFF",X"F7F8FA",X"FEFEFF",X"FCFAFF",X"D28CA4",X"A90C43",X"CA618A",X"F8F5FC",X"FBFFFF",X"FDFDFD",X"FFFFFD",X"FFFFFF",X"F9F8FD",X"FDFDFF",X"FFFFFD",X"FFFEFD",X"FFFDFF",X"FBF1FC",X"AE7178",X"44172B",X"0D0005",X"060709",X"355C6B",X"3A87B3",X"237FB0",X"137D95",X"C3E4F3",X"FFFEFF",X"F5F8EF",X"FBFFFF",X"B9D7FF",X"0396E4",X"00A2DD",X"80B6CE",X"FBFCFF",X"FEFFFF",X"FEFFFF",X"FDFFFC",X"FEFFFF",X"FBFBFD",X"FFF8FF",X"FFFBFF",X"FAFFF9",X"F2F8F6",X"FEFFFF",X"FCFAFB",X"FDFBFC",X"FCFFFF",X"F4FDFC",X"F6FFFA",X"FEF6EB",X"FCFBF9",X"FFFFE6",X"EDE96E",X"D5CF15",X"DAD557",X"F1EFBE",X"E7F1BC",X"E2E0C7",X"DECDC3",X"D3BEC5",X"EED1E3",X"E5BDD7",X"E3C6DC",X"E5BDD8",X"E794BE",X"7D083D",X"38001B",X"64475D",X"FFF0FB",X"FCFFFD",X"F5FFF8",X"FBFBFB",X"FDFAFF",X"FFF5FC",X"FFFEFF",X"86808A",X"120007",X"909599",X"FFF3FF",X"FFF4FF",X"D7F7F2",X"519596",X"0B8F77",X"0E9978",X"306960",X"DDD8DF",X"FFFFFF",X"E8F5EB",X"FFFFF6",X"FBF0B0",X"CDA505",X"E4CC6C",X"F6FFFA",X"F8FFFA",X"FFFDFA",X"FCFCFC",X"FDFEFF",X"FFFCFF",X"FCFDED",X"D1C980",X"A89B00",X"BFB351",X"E8F1DC",X"F8FFFF",X"FFFCFD",X"FEFFFF",X"FBFFFF",X"C7BCC0",X"070004",X"26685A",X"9FD7CE",X"F1FFFF",X"FBFBFD",X"FFFFFB",X"FFFEFD",X"FFFEFD",X"FEFEFC",X"FBFFFC",X"FAFFFC",X"FBFFFC",X"FEFFFA",X"FFFCFD",X"FFFAFC",X"F6EAFE",X"C168B8",X"E216A9",X"CB1A9C",X"FFCAF8",X"F7FFF2",X"FBFEFF",X"FFFBFF",X"D1D2D6",X"041D45",X"16397D",X"C0D5F2",X"FEFFF8",X"FFFBFF",X"FFFFFD",X"FCFCFA",X"FFFFFB",X"FEFDF9",X"FFFDFF",X"FFFAFF",X"FFFCFF",X"C8BCAE",X"19000A",X"BFB0B3",X"FFFDF8",X"FFFEF9",X"FDFCFF",X"FCFCFF",X"FCFBFF",X"FFFEFF",X"E3C7D3",X"7A0500",X"9C110A",X"5F050E",X"5F152E",X"762337",X"4D0304",X"470506",X"A19599",X"FFFCFE"),
(X"FFF8FE",X"FFFAFE",X"BEF3E3",X"1DD599",X"129D73",X"D2D7DA",X"FFFEFF",X"FFEAF7",X"FFCEF3",X"C17CB3",X"7E4E82",X"F9E7FF",X"FFFBF7",X"FFFEF2",X"FFF2FF",X"AF6BA6",X"810073",X"8E018D",X"F0ADF0",X"F1FEEC",X"FEFFF8",X"FFF7FF",X"FFFAFF",X"F9FFFF",X"F9FFFA",X"F6F6F4",X"FFFCFF",X"FFFEFF",X"F6FEFF",X"EFF9FA",X"FFFDFF",X"FFF7FF",X"F2FAFD",X"FFFCFF",X"E3FAF4",X"57CDAB",X"16D99F",X"23D09B",X"B5FFE5",X"FEFFF5",X"F7FFFF",X"F6FEFF",X"FAFFFF",X"FCFFFF",X"FCFFFF",X"FBFCFF",X"FAFBFF",X"FEFFFF",X"F5FDFF",X"FFFAFF",X"EDF8FA",X"FFEEC6",X"FC8D22",X"E76608",X"C18676",X"FFFFEA",X"F9FDFC",X"FFFBFF",X"EBFFF4",X"FFFEF4",X"B3C5E9",X"0849BF",X"7391B7",X"E8F8F8",X"FAFFFF",X"FBFEFF",X"FBFEFF",X"FDFDFF",X"FDFDFF",X"FDFEFF",X"FDFFFC",X"FDFFF9",X"FCFFFF",X"FEF9F3",X"FFFCF1",X"AE9AA5",X"6F4960",X"735C66",X"C3B7C3",X"FFE8FF",X"E6D2ED",X"BB93C8",X"660C52",X"EFDEF0",X"FEFDF9",X"FCFFFF",X"FEFFFF",X"FCFBF6",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FDFDFD",X"FFFAFE",X"FDFEF8",X"CCCAA4",X"9B9A3E",X"C1BE89",X"E8EDB7",X"B4B385",X"C5C585",X"A39280",X"C5D0CA",X"F2FAFF",X"FFFEFF",X"FBFFF1",X"F5FDF0",X"E5F1FF",X"6492C3",X"1276D4",X"0657B2",X"8EBCF7",X"F4FEFF",X"FFFBF4",X"FFFEFF",X"FAFBFF",X"FFFAFF",X"FFF9FC",X"FFFBFC",X"FDFFFE",X"FBFFFF",X"FAFAFC",X"FEFFFF",X"FFFDFD",X"FFE2EA",X"7A5253",X"150103",X"050004",X"D1CED5",X"FFFCFF",X"FBFCFF",X"FBFFFF",X"F1F6FA",X"476ABC",X"000522",X"998A87",X"FFF9F7",X"FCFFFF",X"FBFDFC",X"FFFFFA",X"FFFDFF",X"F2FFFF",X"FFFAFE",X"FFF4FA",X"FFFAFF",X"FAF5FC",X"F8FFFF",X"F0FBF3",X"FFFAF3",X"FF7E8E",X"A50018",X"CA263E",X"99000D",X"FFB3B6",X"FFFCFB",X"FFFAFF",X"EFFFF1",X"FDFEFF",X"FEFEFF",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FBFBFD",X"FAFBFD",X"FEFFFF",X"FEFEFF",X"FCFAFF",X"CF89A1",X"A5083F",X"C85F88",X"F7F4FB",X"FBFFFF",X"FEFEFE",X"FEFEFC",X"FFFFFF",X"FFFEFF",X"FFFFFF",X"FDFCFA",X"FEFAF9",X"FFFAFE",X"FCF2FD",X"AD7077",X"1D0004",X"0F0007",X"AFB0B2",X"E1FFFF",X"A9F6FF",X"74D0FF",X"45AFC7",X"D5F6FF",X"F9F7FC",X"FBFEF5",X"FAFFFF",X"B3D1FF",X"0396E4",X"00A5E0",X"6BA1B9",X"F4F5FA",X"FDFEFF",X"FCFEFD",X"FCFEFB",X"FDFFFE",X"FEFEFF",X"FFFCFF",X"FFFAFF",X"FCFFFB",X"FBFFFF",X"F8F9FB",X"FFFEFF",X"FFFDFE",X"F2F6F7",X"F9FFFF",X"F7FFFB",X"FFFEF3",X"FEFDFB",X"FFFBE0",X"CECA4F",X"D0CA10",X"E8E365",X"FFFECD",X"FEFFD3",X"FFFFE8",X"FFF4EA",X"FFF8FF",X"FFF1FF",X"FFEDFF",X"FFECFF",X"FFF0FF",X"FFB5DF",X"7E093E",X"5B1B3E",X"74576D",X"FFEFFA",X"FCFFFD",X"F1FCF4",X"FFFFFF",X"FFFCFF",X"FFF8FF",X"FAF9FF",X"807A84",X"17000C",X"92979B",X"FFF1FF",X"FFF6FF",X"E3FFFE",X"B3F7F8",X"1DA189",X"1EA988",X"043D34",X"4D484F",X"E2E2E2",X"F7FFFA",X"FBFDF2",X"F7ECAC",X"D1A909",X"E5CD6D",X"F5FFF9",X"F7FFF9",X"FFFDFA",X"FCFCFC",X"FDFEFF",X"FFFAFE",X"F8F9E9",X"CCC47B",X"C6B90A",X"BAAE4C",X"F8FFEC",X"F4FEFF",X"FFF8F9",X"F6F7F9",X"FBFFFF",X"CCC1C5",X"080005",X"26685A",X"98D0C7",X"EEFEFE",X"FAFAFC",X"FEFDF9",X"FFFDFC",X"FFFEFD",X"FFFFFD",X"FCFFFD",X"FAFFFC",X"FAFFFB",X"FDFEF9",X"FFFCFD",X"FFF8FA",X"FFF4FF",X"D47BCB",X"C6008D",X"C11092",X"FAC5F3",X"F8FFF3",X"FAFDFF",X"FFF6FB",X"D0D1D5",X"000C34",X"002165",X"B6CBE8",X"FBFEF5",X"FFF9FF",X"FFFFFD",X"FEFEFC",X"FFFFFB",X"FCFBF7",X"FFFCFF",X"FEF9FF",X"FFFAFF",X"C1B5A7",X"110002",X"BDAEB1",X"FFFFFA",X"FFFFFA",X"F9F8FD",X"FBFBFF",X"FEFDFF",X"FFFEFF",X"E9CDD9",X"6B0000",X"8A0000",X"FFA9B2",X"FFD4ED",X"FFCDE1",X"FFB6B7",X"611F20",X"908488",X"FFFDFF"),
(X"F4FEFD",X"F9FFFF",X"B4EDDC",X"00DB91",X"00D790",X"C0FFEE",X"F0FFFF",X"EBFFFF",X"FEFEFF",X"EFDCF0",X"B2A7B7",X"FDFEFF",X"FCFBF6",X"FCFFFB",X"F7F7FF",X"8F7696",X"5F1262",X"6B017D",X"E4AFF7",X"EBFFF0",X"F0FFEC",X"FFFEFC",X"FFFCFF",X"FFF4FF",X"F5FFFF",X"FAFCFF",X"FDF7FF",X"FFFCFF",X"FBFCFE",X"FBFFFA",X"FEFFFD",X"FFFCFD",X"F5FFFD",X"F8FAF9",X"D1FDF0",X"43D4AB",X"03E2A1",X"07D499",X"9CFFE8",X"F4FFFA",X"FDF7FF",X"FFFDFF",X"FFF9FF",X"FEF7FE",X"FFFCFF",X"FCFAFD",X"FFFFFF",X"FEFFFD",X"FCFCF2",X"FFFBFF",X"FCFFFF",X"FFDBB8",X"F57D0C",X"DB7200",X"9F7E6B",X"FFFEFF",X"FFFFF6",X"FFF7FE",X"EDFFFA",X"FFFFF0",X"B5D8EE",X"004EBE",X"6997C8",X"E3F5FF",X"FFFAFB",X"FFFAFB",X"FFF8FD",X"FFF9FF",X"FFFAFE",X"FFFFFF",X"FAFFFB",X"F9FFFB",X"FFFEEF",X"FFF7FF",X"FFFAFF",X"AF7AAE",X"630168",X"AA65A6",X"FFF7F8",X"FCFAFF",X"FFFAFF",X"FFF6FF",X"C68EBD",X"EAE7F2",X"FFFCFD",X"FFFDFF",X"FDFDFF",X"FCFDF8",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FDFDFD",X"EFFFF3",X"FFFFE6",X"F7D886",X"E3B70C",X"F5D156",X"F1F2A6",X"F0F4DD",X"FAE9D9",X"FFFCEF",X"FDFEFF",X"F7F6FF",X"FFFDFF",X"FEFFED",X"F6FFEC",X"ECFFFF",X"93BEE8",X"0163C6",X"0465CE",X"64A8F1",X"EAFFFF",X"FBFEF7",X"F9FCFF",X"FAFEFF",X"FFFFEC",X"F1FFFF",X"FFFEFF",X"F6FFFF",X"F8FCFF",X"FFF8FF",X"F1FFFF",X"F0FDFF",X"FFC6E7",X"AC2533",X"66151B",X"130000",X"D3CDCD",X"FFFDFF",X"F7F5FA",X"F8FFFF",X"E2F7FA",X"3F72CB",X"000643",X"8D838E",X"FDF6EE",X"F6FAF9",X"FCFDFF",X"FFFBFF",X"FFFDFA",X"FDFBFE",X"F8FFFF",X"FBFFFF",X"F8FCFD",X"F7FFFF",X"FAFDFF",X"FFF6FB",X"FCFDF8",X"EBB6C6",X"98050F",X"D0161B",X"A93039",X"F6CDDD",X"FFF9FF",X"FFFDFF",X"F7FFFB",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FCFFFF",X"FEFEFF",X"FEFFFD",X"A6858C",X"6D001F",X"C46688",X"FBF6FC",X"F8FFFE",X"FFFBFB",X"FFFFFD",X"FFFFFF",X"FCFCFE",X"FCFCFC",X"FFFFFD",X"FFFEFD",X"FFF9FD",X"FDF3FC",X"9F698B",X"070009",X"726B72",X"FDF4F9",X"F5FFFF",X"EDFFFF",X"E7FFFF",X"B6CFC9",X"ECF8F8",X"F3F7FF",X"F5FEFF",X"FFFFF6",X"BBDFED",X"00A3DD",X"00A8EC",X"648AB7",X"F6F5FA",X"FDFEFF",X"FBFCFE",X"FFFFFF",X"FDFBFC",X"FDF7FB",X"FFFCFF",X"FFFBFF",X"FAFFFF",X"FFFFFD",X"FDF8F5",X"FFFAFB",X"FDF7F7",X"FFFEFB",X"F5F6F1",X"F9FFFF",X"FFFCFF",X"F9FEFF",X"FCFEF1",X"DAD255",X"D1D200",X"DFE672",X"FBFCFF",X"FDFDF1",X"F5FFF8",X"FBFBF9",X"F9FBFA",X"FAF9F7",X"FEF6F4",X"F3F9F7",X"FDFBFF",X"F0C5E3",X"B8004D",X"C10B60",X"B74580",X"FFEAFF",X"FFFEFF",X"F8FAF5",X"F6FBF7",X"FFFDFF",X"F3FFFF",X"FDF0FF",X"C36D9A",X"92003D",X"D6A6BE",X"FFF1FA",X"FBFCFF",X"F1FFFF",X"F7FFFF",X"B5E2DB",X"4F8D80",X"31564F",X"000807",X"595758",X"F4F2F3",X"FFFDFF",X"F7EFC0",X"A88B13",X"E2CE89",X"FCFFFF",X"F6F7F1",X"FFFCF6",X"FFFDFF",X"FAFFFF",X"F9FFFB",X"FFFAEA",X"DAC087",X"B79C00",X"DAC15A",X"FAF4DE",X"F8FBFF",X"FAFDF2",X"FFF9FF",X"FFFBFA",X"CFC5C6",X"000602",X"01332A",X"72CBB7",X"DAFFFE",X"FFF8FF",X"FFFCFF",X"FFFCFF",X"FFFAFF",X"FEF9FF",X"FFFEFF",X"FEFFFF",X"FDFAFF",X"FFFCFF",X"FFFBF9",X"FFF9FB",X"F7E6F9",X"D479C9",X"E01AAD",X"B3088C",X"FFC9FA",X"FCFFF2",X"F8FDFF",X"FFFDFF",X"CCC8BF",X"00020E",X"000732",X"BAC6DE",X"FAFDF6",X"FFFDFF",X"F8FEFC",X"FFFFF8",X"FFFAF4",X"FFFCFF",X"FFFCFF",X"F4F7FC",X"F1FFFF",X"8CA9C7",X"00013C",X"ADB4D0",X"FFFDF7",X"FCFDEF",X"F8FFFF",X"F7FFFF",X"F9F7FF",X"FFFAFF",X"D1D3D0",X"100005",X"665355",X"ECEEEB",X"FEFFFF",X"FFFBFF",X"FFFAFF",X"D9CED6",X"CFC7C4",X"FFFFFA"),
(X"F5FFFE",X"F6FFFE",X"BCF5E4",X"00DD93",X"03E39C",X"AFEEDD",X"EFFFFF",X"EAFFFF",X"F5F5FF",X"FFF7FF",X"F6EBFB",X"FEFFFF",X"F8F7F2",X"FBFFFA",X"FCFCFF",X"947B9B",X"510454",X"650077",X"E2ADF5",X"F1FFF6",X"EEFFEA",X"F6F5F3",X"FFFCFF",X"FFF5FF",X"F0FEFF",X"FBFDFF",X"FFFCFF",X"FFFBFF",X"F8F9FB",X"FCFFFB",X"FEFFFD",X"FDF9FA",X"F3FFFB",X"FEFFFF",X"D9FFF8",X"47D8AF",X"05E4A3",X"0BD89D",X"8BF7D7",X"EEFBF4",X"FFFAFF",X"FCF7FE",X"FFFCFF",X"FDF6FD",X"FEF7FE",X"FFFEFF",X"F8F8F8",X"FEFFFD",X"FFFFF6",X"FFFBFF",X"F5F9FA",X"F6CEAB",X"EC7403",X"E77E08",X"C7A693",X"FAF9FF",X"FDFDF3",X"FFF9FF",X"F1FFFE",X"FCFAEB",X"ACCFE5",X"0660D0",X"5A88B9",X"DFF1FF",X"FFF6F7",X"FFF8F9",X"FFFAFF",X"FFF5FB",X"FFFDFF",X"F7F7F7",X"F6FBF7",X"F9FFFB",X"FFFEEF",X"FFF7FF",X"FDF4FF",X"B37EB2",X"630168",X"A762A3",X"F8EEEF",X"FCFAFF",X"FFFAFF",X"FFF4FF",X"FFD6FF",X"FFFDFF",X"FFF6F7",X"FFFDFF",X"FFFFFF",X"FFFFFB",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FDFDFD",X"E8FDEC",X"FFFFE3",X"ECCD7B",X"D3A700",X"E3BF44",X"FEFFB3",X"F4F8E1",X"FFFCEC",X"FFFBEE",X"FDFEFF",X"FAF9FF",X"FFFEFF",X"FEFFED",X"F8FFEE",X"EEFFFF",X"A5D0FA",X"005BBE",X"0B6CD5",X"5B9FE8",X"E0F8FF",X"FEFFFA",X"F9FCFF",X"FBFFFF",X"FFFFED",X"F5FFFF",X"FFFEFF",X"F8FFFF",X"FBFFFF",X"FFF6FF",X"EAFDFF",X"F5FFFF",X"F0ADCE",X"910A18",X"611016",X"5D4342",X"F6F0F0",X"FFFDFF",X"FFFEFF",X"F8FFFF",X"E2F7FA",X"4376CF",X"000340",X"796F7A",X"FFFCF4",X"FCFFFF",X"FBFCFF",X"FFFDFF",X"FDF9F6",X"FDFBFE",X"F8FFFF",X"F5FBF9",X"FBFFFF",X"F4FFFF",X"F4F7FC",X"FFFCFF",X"FFFFFB",X"FFCADA",X"C4313B",X"B90004",X"CE555E",X"FFEBFB",X"FFF7FF",X"FFFDFF",X"F3FFF7",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FCFFFF",X"FCFCFE",X"F4F6F3",X"AA8990",X"5B000D",X"BA5C7E",X"F6F1F7",X"F9FFFF",X"FFFCFC",X"F9F9F7",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFD",X"FFFDFC",X"FFFAFE",X"FFF5FE",X"945E80",X"0C000E",X"807980",X"FFFAFF",X"F2FCFE",X"ECFFFF",X"E9FFFF",X"EDFFFF",X"F2FEFE",X"F6FAFF",X"F8FFFF",X"FFFFF6",X"BFE3F1",X"0096D0",X"00B1F5",X"557BA8",X"F2F1F6",X"FEFFFF",X"FEFFFF",X"F1F1F1",X"FFFEFF",X"FFFDFF",X"FAF3FB",X"FFFBFF",X"F8FEFE",X"FAFAF8",X"FFFEFB",X"FFFCFD",X"FFFDFD",X"FDF8F5",X"FFFFFB",X"F7FFFF",X"FFFCFF",X"F3F8FE",X"FFFFF4",X"E7DF62",X"DCDD06",X"D6DD69",X"F6F7FB",X"FFFFF4",X"F5FFF8",X"FEFEFC",X"FCFEFD",X"FFFEFC",X"FFFDFB",X"FBFFFF",X"FFFDFF",X"EEC3E1",X"BD0052",X"B90358",X"BC4A85",X"FFE0F5",X"FFFEFF",X"FEFFFB",X"FAFFFB",X"FFFCFF",X"F5FFFF",X"F2E5F6",X"BC6693",X"A30E4E",X"DFAFC7",X"FFF8FF",X"FCFDFF",X"EFFFFF",X"EFFAFC",X"DDFFFF",X"A7E5D8",X"41665F",X"161F1E",X"060405",X"706E6F",X"FAF4F8",X"FFF9CA",X"A88B13",X"D4C07B",X"F7FBFC",X"FFFFFA",X"FFF9F3",X"FFFDFF",X"F9FEFF",X"F3FDF5",X"FFFBEB",X"D8BE85",X"BDA200",X"C1A841",X"F9F3DD",X"FCFFFF",X"FEFFF6",X"FFF8FF",X"FFFEFD",X"CEC4C5",X"000804",X"1C4E45",X"62BBA7",X"D8FFFC",X"FFF4FE",X"FFFAFF",X"FFFCFF",X"FFF8FF",X"FFFDFF",X"F8F7FD",X"FBFCFF",X"FFFDFF",X"FFF8FF",X"FFF7F5",X"FFF4F6",X"FFF4FF",X"B055A5",X"C1008E",X"FF55D9",X"FFD0FF",X"FEFFF4",X"EFF4F8",X"FCF6F8",X"D4D0C7",X"000410",X"00042F",X"A4B0C8",X"FEFFFA",X"FFFBFF",X"FBFFFF",X"F4F5ED",X"FFFEF8",X"FFFCFF",X"FEF7FE",X"FCFFFF",X"E5F7FF",X"829FBD",X"00114C",X"B9C0DC",X"FFFEF8",X"FFFFF3",X"F4FEFF",X"F7FFFF",X"FDFBFF",X"FFF6FB",X"CCCECB",X"100005",X"6F5C5E",X"E8EAE7",X"FBFCFF",X"FCF7FD",X"FFFDFF",X"FFF7FF",X"FDF5F2",X"FCFBF6"),
(X"F8FFFF",X"ECFFFD",X"A3EBD5",X"12DA99",X"00D08E",X"9FEDD7",X"EEFAFA",X"FFFEFF",X"FFF4FF",X"FFF5FD",X"FAFBF5",X"F8FFFA",X"FFFEFD",X"F7F2F8",X"FAFDFF",X"CFC5D0",X"0A000C",X"5B0860",X"B952BD",X"FFD5FF",X"FFEFFF",X"FEFDFF",X"FBFFFB",X"FBFFF7",X"FFFBFF",X"FDFDFD",X"FAFFFE",X"FAFAF8",X"FFFBF5",X"FBFBF3",X"EFFFF8",X"E6FFFF",X"EAFFF3",X"FEFFFD",X"F8FFFF",X"AFEFE1",X"28BF96",X"04D699",X"3FE9BA",X"C0FFF8",X"FEFFFF",X"FAF8F9",X"F8F4F5",X"FFFDFF",X"FFFCFC",X"FEFDF9",X"FEFFFA",X"F8FEF4",X"F5EFE3",X"FFFCF8",X"FFFBE1",X"FCB76A",X"F47E02",X"D78829",X"F8EDD9",X"FBFFFF",X"F9F8FD",X"FFF8FF",X"F7FBFC",X"FFFFF8",X"9AC6EB",X"0765C5",X"3B6DA0",X"DADDFE",X"F8FFFD",X"F3FCF7",X"FCFFFB",X"FCFDF8",X"FFFFFB",X"FDFCF8",X"FFFFFD",X"FFFFFD",X"FCFCFF",X"F5F5FD",X"FFF5FF",X"B56DB6",X"78077B",X"A964B4",X"FAFBF6",X"F8FFF9",X"F6FFEC",X"EEFFFA",X"F8FFFF",X"FAFEFF",X"FFF1FC",X"FFF9FB",X"FEFAF9",X"F7FCFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FDFDFD",X"F7FFED",X"FFFBE8",X"E2CB7F",X"DAB21F",X"ECBD51",X"FFF9C5",X"F9FFFB",X"FBEFFB",X"FCFDFF",X"FDFEFF",X"FFFEFF",X"FFFCFA",X"FFFEF8",X"FFFDFC",X"F7FEFF",X"D4E6F4",X"1967BC",X"147BF1",X"0661CC",X"AADEFF",X"EEFFF6",X"FEFFF6",X"FDF4F7",X"FDF8F2",X"EBFFF6",X"FFF9F9",X"F9F5F4",X"FCFDF8",X"FFFFFA",X"E8FDEE",X"FFFAF6",X"FF8BA8",X"B8000B",X"890016",X"CC95A8",X"F9FFFF",X"F9FFF8",X"FFF5EF",X"FEFBFF",X"D3EEFF",X"2066C5",X"001F79",X"616884",X"EDF3F1",X"F8FDFF",X"F2F3F8",X"F7F7FF",X"F8FFFF",X"FFF6FF",X"F1F7F5",X"F7FDF9",X"FAF8F9",X"FBFFFF",X"FFF7FF",X"FFF4FF",X"FDF2F6",X"FFE3F2",X"B85E55",X"BE0007",X"E07684",X"FBFCFF",X"FAF5F9",X"FAFCFB",X"FFF8FF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FFFFFD",X"F6FBF7",X"817778",X"5C001D",X"C04F7B",X"FEE2F1",X"FEFFFF",X"FFFAF8",X"FFFFFD",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FDFEF9",X"FAF9F5",X"FFFAFE",X"F7F0F8",X"6C5F56",X"000B0A",X"739A97",X"EBFFF7",X"FDFAF3",X"FFFBFF",X"F0F9FF",X"FFF6FC",X"FFFDF4",X"FFFCF6",X"F3F5F2",X"FDF8F2",X"EFFDFE",X"57BBDD",X"15A0DB",X"045A95",X"AAB3BA",X"F4FFFF",X"F1FCFF",X"F9FFFF",X"F7FAF1",X"F3F5EA",X"FBFFFB",X"F4FEFD",X"FFFDFF",X"FFF7F8",X"FFFDFF",X"F8FCFF",X"F7FBFF",X"FFFCFF",X"FAEEEE",X"FFFBFF",X"FFFBFF",X"F6FDF5",X"FFFFDF",X"EADD53",X"DAD600",X"DEE564",X"FCFEFD",X"FFFEFF",X"F6FFF9",X"FFFFFB",X"FEFFFA",X"FFFFF5",X"FFF9F5",X"F8F6F7",X"FFF5FF",X"FBBDEC",X"8C0842",X"B31359",X"B6477C",X"FFECFF",X"FCF7FB",X"FEFAF7",X"FBFFFC",X"FAFAFA",X"FAF2FD",X"FFDBFD",X"DA5199",X"BA0055",X"E8B1D0",X"F8FFFF",X"F4F8F9",X"FFF4FF",X"F8FFFA",X"FBFFFD",X"F3FDFE",X"BAC8C8",X"000604",X"221E1F",X"090A0F",X"758489",X"C1D1C4",X"000700",X"A29E95",X"FFFDFF",X"F9F6EF",X"FFFAFF",X"FBF3FF",X"F8FFF3",X"F7FFF8",X"F4EDE3",X"C2A98B",X"C2AD2E",X"AE9D27",X"FEEFD0",X"FFFEFF",X"F5FFF3",X"FEFFFF",X"F5FBF7",X"ECEBE9",X"29423C",X"254240",X"46A891",X"AEF5E7",X"FBFFFF",X"F9FFFD",X"F6FBF7",X"F4F6F1",X"FCFFF8",X"F5FCF4",X"F9FFF9",X"FBFBF9",X"FFFDFD",X"FFFFFB",X"F3F5FF",X"FFCAFF",X"E74AB3",X"A10E76",X"DCA0DC",X"FBF8FF",X"FAF8FD",X"FCFFFF",X"FFFFFD",X"D9D5CA",X"434343",X"020318",X"A1A0B2",X"FFFEFF",X"F9F5F2",X"F7FFFF",X"FEFCFD",X"FFFBFF",X"FBF5F7",X"FFFFEE",X"F1FAE9",X"DBF6FF",X"5D88E4",X"00287E",X"B0BEEB",X"FEF8FA",X"FFFFF5",X"ECFBF6",X"F5FFFF",X"FBFBF9",X"FFFDF8",X"B7D1E2",X"000D6A",X"546AC0",X"EDE9FF",X"FFF7FD",X"FFF7F6",X"F2F8FF",X"F3F8FC",X"FFFFFF",X"F9FFFF"),
(X"F9FFFF",X"E9FFFA",X"A5EDD7",X"06CE8D",X"04D593",X"93E1CB",X"F4FFFF",X"FDFBFF",X"FFF4FF",X"FFF7FF",X"FEFFF9",X"F1FDF3",X"FEFAF9",X"FFFDFF",X"FCFFFF",X"FEF4FF",X"6E5D70",X"5D0A62",X"630067",X"CF91D0",X"FFEEFF",X"F9F8FD",X"F7FEF7",X"F6FCF2",X"FDF2F6",X"F9F9F9",X"FBFFFF",X"FFFFFD",X"FFFEF8",X"F9F9F1",X"EFFFF8",X"CFF5EA",X"E5FBEE",X"F6F8F5",X"F8FFFF",X"BEFEF0",X"42D9B0",X"12E4A7",X"13BD8E",X"B4FDEC",X"FAFCFB",X"FEFCFD",X"FFFEFF",X"FFFDFF",X"FCF6F6",X"FDFCF8",X"F7FAF3",X"FCFFF8",X"FFFFF3",X"FFFCF8",X"F4E3C9",X"D59043",X"EF7900",X"F2A344",X"F8EDD9",X"FBFFFF",X"FAF9FE",X"FFF9FF",X"F4F8F9",X"FFFFF7",X"8EBADF",X"0664C4",X"023467",X"D6D9FA",X"F8FFFD",X"F3FCF7",X"FCFFFB",X"FDFEF9",X"F7F6F2",X"FFFFFB",X"FEFEFC",X"FEFEFC",X"FEFEFF",X"FBFBFF",X"FFF0FF",X"9F57A0",X"710074",X"A762B2",X"FAFBF6",X"F6FFF7",X"FBFFF1",X"E8FFF4",X"EFF9FA",X"F3F7FF",X"FFF6FF",X"FFF9FB",X"FCF8F7",X"FBFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FDFDFD",X"F3FFE9",X"FFFFEC",X"E8D185",X"D9B11E",X"EABB4F",X"FEF2BE",X"F6FFF8",X"FFF6FF",X"FCFDFF",X"FCFDFF",X"FFFEFF",X"FFFAF8",X"FFFDF7",X"FFFEFD",X"F7FEFF",X"E8FAFF",X"64B2FF",X"076EE4",X"0863CE",X"71A5CC",X"E5FDED",X"FDFFF5",X"FFFCFF",X"FFFEF8",X"EBFFF6",X"FFFDFD",X"FFFEFD",X"FFFFFB",X"FAFBF5",X"EEFFF4",X"FFF1ED",X"E16683",X"B60009",X"990F26",X"FFDCEF",X"F9FFFF",X"EAF4E9",X"FFFCF6",X"FFFDFF",X"C7E2F5",X"1A60BF",X"1B3A94",X"444B67",X"DFE5E3",X"FBFFFF",X"FEFFFF",X"F8F8FF",X"F9FFFF",X"FFECF9",X"FBFFFF",X"FBFFFD",X"FDFBFC",X"FAFFFF",X"FFF9FF",X"FFF4FF",X"FFFBFF",X"FFF2FF",X"C1675E",X"BA0003",X"E77D8B",X"EFF0F5",X"FFFDFF",X"FEFFFF",X"FFF8FF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FDFFFE",X"FDFFFE",X"FDFFFE",X"FCFBF9",X"FAFFFB",X"7C7273",X"5E001F",X"BB4A76",X"FEE2F1",X"FEFFFF",X"FEF6F4",X"FFFFFD",X"FEFEFE",X"FAFAFC",X"FCFCFC",X"FEFFFA",X"FDFCF8",X"FFFDFF",X"F0E9F1",X"5F5249",X"000807",X"85ACA9",X"E8FFF4",X"FCF9F2",X"FCF4FF",X"F8FFFF",X"FFF9FF",X"FFFCF3",X"FFFBF5",X"FEFFFD",X"FEF9F3",X"F3FFFF",X"82E6FF",X"0691CC",X"095F9A",X"000209",X"D1DCE2",X"F5FFFF",X"F5FEFB",X"FBFEF5",X"FFFFF6",X"FBFFFB",X"F1FBFA",X"FFFDFF",X"FFF6F7",X"F8F2F4",X"FBFFFF",X"E2E6EF",X"DFD6D9",X"FFF9F9",X"FFFCFF",X"FFFAFE",X"FBFFFA",X"FCFCDA",X"EADD53",X"D8D400",X"EBF271",X"FEFFFF",X"FEFCFF",X"F6FFF9",X"FFFFFB",X"FAFDF6",X"FFFFF5",X"FFFCF8",X"FBF9FA",X"FFF8FF",X"FEC0EF",X"720028",X"96003C",X"A13267",X"FFE6FA",X"FFFAFE",X"FFFBF8",X"FBFFFC",X"FEFEFE",X"FFFAFF",X"FFD6F8",X"C23981",X"B60051",X"F4BDDC",X"F9FFFF",X"FCFFFF",X"FFF5FF",X"F2FEF4",X"F2F8F4",X"F6FFFF",X"F5FFFF",X"A2A8A6",X"030000",X"232429",X"000409",X"334336",X"040E00",X"949087",X"FDF8FE",X"FFFFF8",X"FFFAFF",X"FFFBFF",X"EEFBE9",X"F3FFF4",X"F8F1E7",X"72593B",X"B7A223",X"CAB943",X"FBECCD",X"FFFEFF",X"F0FCEE",X"FCFDFF",X"FBFFFD",X"FFFFFD",X"839C96",X"000907",X"3EA089",X"86CDBF",X"F4F9FD",X"F4FDF8",X"F6FBF7",X"FEFFFB",X"F4F7F0",X"F4FBF3",X"FBFFFB",X"F9F9F7",X"FFF9F9",X"F4F5F0",X"F9FBFF",X"F7B3EC",X"D2359E",X"C8359D",X"FFCBFF",X"FFFCFF",X"F9F7FC",X"F5F9FC",X"FFFEFC",X"FEFAEF",X"3A3A3A",X"000013",X"A3A2B4",X"FFFDFE",X"FCF8F5",X"F5FFFE",X"F8F6F7",X"FFF5FD",X"FFFDFF",X"F6F7E5",X"FBFFF3",X"D7F2FF",X"345FBB",X"1C4AA0",X"C2D0FD",X"FFF9FB",X"FFFFF6",X"F1FFFB",X"F7FFFF",X"FAFAF8",X"FFFDF8",X"ABC5D6",X"0B2582",X"5369BF",X"EBE7FF",X"FFF5FB",X"FFF8F7",X"F4FAFF",X"FBFFFF",X"F0F0F2",X"FBFFFF"),
(X"FFF9FE",X"F5F9FA",X"8BF3D2",X"00D78B",X"00D993",X"7FE2C5",X"E9FFFE",X"F2FAFC",X"FCFBFF",X"F4FFFE",X"DDFFF8",X"CBFAE8",X"F7FDFD",X"FFF4FB",X"FBF2F5",X"FFFAFD",X"D4CCC9",X"39022C",X"9C2C92",X"70006B",X"D586D7",X"FFDCFF",X"FFEEFF",X"FEFCFD",X"FFF4FF",X"FFFAFF",X"FFF2F9",X"FFEFF4",X"FFF8F8",X"F5FFFD",X"C8FFFC",X"4FBAA6",X"BBE6D5",X"F7FFFF",X"FBFAFF",X"E9FBFB",X"91E5CD",X"19C690",X"36EEB8",X"3EB99A",X"D4EBE3",X"F2FFFF",X"EEF8FA",X"F7F7FF",X"FFFDFF",X"FFFDFF",X"F8F8FF",X"F7FBFF",X"FFF4FF",X"FFF9FA",X"AA917B",X"C48C42",X"C98436",X"F7D2B5",X"FFFFF6",X"FDFFF2",X"FFFAFF",X"FFFDFF",X"FEFDFF",X"F0EFEB",X"8597BD",X"1E4767",X"000204",X"FBD6C6",X"FEFEFF",X"FFFCFF",X"FFFDFF",X"FFF9F6",X"FFFDF8",X"F5EEE8",X"EDE8E5",X"FFFEFD",X"F2F7FD",X"F4FFEE",X"D8E8DE",X"5D4553",X"38002F",X"8D7396",X"F6F7E7",X"FFEFEE",X"FFF9FF",X"FBF2F5",X"FEFDFF",X"FFD5FF",X"FFE3FF",X"FFFEFB",X"FCFFF6",X"FFFBFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FDFDFD",X"FFF7F7",X"FFE7F4",X"959070",X"4B4A12",X"BBA677",X"FCF0D8",X"F5FFE9",X"FBFFFF",X"FBFEFF",X"FDFDFD",X"FFFFFB",X"FFFBFA",X"FFF9FE",X"FFFCFF",X"FCFBFF",X"FFFFFF",X"D0ECF0",X"165C98",X"2679F1",X"1561D9",X"7DC8FF",X"DBFFFF",X"F2F9FF",X"F7F7F5",X"FFF6FF",X"FFEEFC",X"FFF8FF",X"F7FEF7",X"F2FDED",X"FFF6ED",X"FFA5AC",X"A3071C",X"8B030F",X"F7ADBA",X"F9E9F6",X"FCF9FF",X"FFFEF8",X"FCFEF3",X"F7FEFF",X"C4C8E5",X"165BB8",X"183B95",X"0B1A31",X"E4E7EC",X"FFF9FF",X"FFEFE2",X"FFF8F3",X"F3F8FC",X"FFF8FF",X"F1E2E7",X"EEDEDF",X"FFFAFB",X"FFF7FD",X"FFFCFF",X"FFFBFF",X"FCFFFF",X"FFE7EF",X"D75A62",X"C8000C",X"DB6170",X"FBEFEF",X"F9F4F1",X"FFFEFD",X"FDFAFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FDFFFE",X"FDFFFE",X"FEFEFE",X"FEFEFE",X"FDFDFD",X"E2E6E5",X"59545A",X"68002B",X"CE3176",X"FFC3E9",X"FFF6FF",X"FFFEFD",X"FFFEFC",X"FCFCFC",X"FDFDFF",X"FEFFFF",X"FEFFFB",X"FBFCF7",X"FFFEFF",X"DBD8DF",X"433245",X"00224B",X"79AEE2",X"EDFFFF",X"F5FFF8",X"FDEEFF",X"FFF4FF",X"F4FAEE",X"FFF6F9",X"F5EDDA",X"FCFCF4",X"F9F7FF",X"FFFDFF",X"ECF6FF",X"6BA8C7",X"238FB5",X"003F5F",X"0C4E6E",X"A4D7F6",X"E9FFFF",X"F2F8FF",X"FFF5FD",X"FFFAFF",X"FFFBFF",X"FAF5FB",X"FEFFFF",X"E7FFFF",X"CFFFFF",X"6093AE",X"314550",X"FFFDFF",X"FFF5F9",X"F9FCFF",X"FFFAEE",X"FFF4B6",X"EBDA46",X"E3D80D",X"EAE34C",X"FFFDCA",X"FAF9FF",X"FFFAFF",X"FFF9FF",X"F7F4FF",X"FEFFFF",X"FFFFFA",X"F2FFF3",X"F9FFF5",X"D8B3BB",X"000300",X"150000",X"49202E",X"D7CCD2",X"F9FFFF",X"FCFFFD",X"FBF9FA",X"FFFAFE",X"F9FFFF",X"F9BFE7",X"B10D66",X"C3005D",X"F6A3D1",X"F5F3F8",X"F8FFFF",X"FFFBFF",X"FFFBF8",X"FFFCFE",X"F6F9FE",X"F3F6FB",X"FBFFFF",X"A7B8B2",X"13423A",X"2E776C",X"20615B",X"003034",X"789AA6",X"FFFDFF",X"FCFBF6",X"FAF4FF",X"FFF5FF",X"F7FFEF",X"FFFFFD",X"F2F7F1",X"555648",X"AFAF57",X"AFB223",X"F8F5C0",X"FFFFFD",X"FCFFFD",X"F7FFFF",X"F3FCF7",X"FAFBF6",X"E2E0E1",X"323A3D",X"3B6460",X"456F6B",X"B2C4C6",X"FBFFFF",X"FAFBFF",X"FCFAFD",X"FFFDFF",X"FEFCFF",X"FFFCFF",X"FFF2FB",X"FFF3FF",X"FFF2FF",X"FFD2FF",X"E056B5",X"A71874",X"EBADDE",X"FFF7FF",X"FEFDFF",X"F2FFFF",X"FEFDFF",X"F9FBF8",X"FCFCFC",X"8E8389",X"0F0006",X"514354",X"E5DDEC",X"FDFEF9",X"F6FBFE",X"FFFCFF",X"FFFAFF",X"F9FFFF",X"FBFFFA",X"FCFFFF",X"CEDEFF",X"12388D",X"6182B5",X"E7F2FF",X"FFFEFF",X"FBFBF9",X"F8FCFB",X"FFFFFA",X"F8F8F6",X"F2FDFF",X"9CB8E7",X"063FB0",X"1C5FB8",X"C5E6FF",X"F7FEFF",X"F9FFEF",X"F2FBF6",X"FEFAFB",X"F1FCFF",X"EEFFFF"),
(X"FFF8FD",X"F9FDFE",X"79E1C0",X"00DF93",X"00D690",X"82E5C8",X"E0F9F5",X"F7FFFF",X"FAF9FE",X"F7FFFF",X"D0FCEB",X"97C6B4",X"E7EDED",X"FFFAFF",X"FFFCFF",X"FDEEF1",X"FEF6F3",X"D69FC9",X"66005C",X"8D1488",X"641566",X"AD81B2",X"F5DEFA",X"FEFCFD",X"FFF4FF",X"FFFAFF",X"FFFAFF",X"FFF8FD",X"FFFAFA",X"F1FFF9",X"B4F6E8",X"38A38F",X"C6F1E0",X"EFFBF9",X"FCFBFF",X"F2FFFF",X"C2FFFE",X"3AE7B1",X"12CA94",X"0C8768",X"2C433B",X"D1E4E0",X"F8FFFF",X"F9F9FF",X"FFFDFF",X"FCFAFF",X"FEFEFF",X"FBFFFF",X"FFF9FF",X"A3999A",X"160000",X"9F671D",X"FFC375",X"FFF7DA",X"F9F9EF",X"FCFFF1",X"FFFBFF",X"F9F6FD",X"FFFEFF",X"FFFFFB",X"596B91",X"000D2D",X"000507",X"E5C0B0",X"FEFEFF",X"FFFCFF",X"FFFDFF",X"FFF8F5",X"F9F0EB",X"7B746E",X"A39E9B",X"FFFBFA",X"F5FAFF",X"F5FFEF",X"CBDBD1",X"14000A",X"220019",X"82688B",X"FFFFF1",X"FFF6F5",X"FFF7FF",X"FFFCFF",X"F7F6FF",X"95699A",X"D2B0D5",X"FFFCF9",X"FCFFF6",X"FDF7FF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FDFDFD",X"FFFBFB",X"EED6E3",X"130E00",X"080700",X"685324",X"F5E9D1",X"F9FFED",X"EAEFF2",X"FBFEFF",X"FDFDFD",X"FCFDF8",X"FFFDFC",X"FFF8FD",X"FFFCFF",X"FCFBFF",X"FFFFFF",X"DEFAFE",X"9AE0FF",X"085BD3",X"1864DC",X"216CAF",X"A5D1EA",X"EEF5FD",X"FFFFFD",X"FFF8FF",X"FFF7FF",X"FFFBFF",X"F9FFF9",X"F8FFF3",X"F0CFC6",X"B64D54",X"95000E",X"FD7581",X"FFE0ED",X"FFF9FF",X"FDFAFF",X"FFFBF5",X"FFFFF6",X"F7FEFF",X"B3B7D4",X"0D52AF",X"2D50AA",X"00041B",X"DDE0E5",X"FFFBFF",X"FFEFE2",X"FFFDF8",X"FBFFFF",X"FAE6F1",X"594A4F",X"C0B0B1",X"FFFAFB",X"FFFBFF",X"FFF9FF",X"FFFAFE",X"F7FBFA",X"F8DAE2",X"C64951",X"CF0013",X"C24857",X"EEE2E2",X"FFFEFB",X"F7F3F2",X"FFFDFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FDFFFE",X"FDFFFE",X"FDFFFE",X"FEFEFE",X"FDFDFD",X"FFFFFF",X"DFE3E2",X"050006",X"8C214F",X"AB0E53",X"FFB7DD",X"FAF0F9",X"FFFDFC",X"FFFFFD",X"FFFFFF",X"FFFFFF",X"FDFFFE",X"FAFCF7",X"F8F9F4",X"FFFEFF",X"CFCCD3",X"0C000E",X"115A83",X"84B9ED",X"ECFFFF",X"F2FFF5",X"FFF8FF",X"FFF7FF",X"FCFFF6",X"BBACAF",X"D2CAB7",X"FFFFF8",X"FFFDFF",X"F6F0F2",X"F7FFFF",X"BAF7FF",X"329EC4",X"347B9B",X"3B7D9D",X"5083A2",X"C9E5FB",X"F8FEFF",X"FFFBFF",X"FEF2FC",X"FFF9FF",X"FFFCFF",X"F9FAFE",X"E5FFFF",X"BAF0FF",X"2C5F7A",X"96AAB5",X"FDF7F9",X"FFF6FA",X"F9FCFF",X"FFFBEF",X"FFF4B6",X"D9C834",X"E5DA0F",X"DDD63F",X"FFFECB",X"FFFEFF",X"FFFAFF",X"FFF9FF",X"FCF9FF",X"FEFFFF",X"FBFCF6",X"F1FFF2",X"F9FFF5",X"C29DA5",X"030700",X"36181A",X"2D0412",X"D7CCD2",X"F9FFFF",X"F9FEFA",X"FFFDFE",X"FCF7FB",X"F9FFFF",X"FFC7EF",X"AB0760",X"C5005F",X"E28FBD",X"FFFEFF",X"F3FEFA",X"FFFAFE",X"FFFBF8",X"FEF8FA",X"F5F8FD",X"FCFFFF",X"FBFFFF",X"EAFBF5",X"99C8C0",X"2F786D",X"4F908A",X"307E82",X"93B5C1",X"FFFDFF",X"FFFFFA",X"FFFCFF",X"FFF9FF",X"F1FFE9",X"FFFFFD",X"EDF2EC",X"444537",X"9A9A42",X"999C0D",X"F5F2BD",X"FAF9F7",X"FAFFFB",X"F0FCFA",X"F9FFFD",X"FFFFFB",X"FEFCFD",X"C4CCCF",X"000F0B",X"000D09",X"011315",X"ABB0B4",X"FBFCFF",X"F7F5F8",X"FFFEFF",X"FFFEFF",X"FFFDFF",X"FFF6FF",X"FFF7FF",X"F0D2F6",X"C27EBB",X"B22887",X"FF8AE6",X"FFD7FF",X"FFFBFF",X"F7F6FB",X"F3FFFF",X"FFFEFF",X"F6F8F5",X"FFFFFF",X"D1C6CC",X"190810",X"08000B",X"857D8C",X"EFF0EB",X"F4F9FC",X"FFFCFF",X"FFFAFF",X"EEF4F4",X"FBFFFA",X"EFF2F9",X"7787BA",X"00166B",X"ABCCFF",X"F4FFFF",X"FCF8F9",X"F7F7F5",X"F9FDFC",X"FAF9F4",X"FDFDFB",X"F7FFFF",X"7A96C5",X"0D46B7",X"1356AF",X"B5D6FF",X"EFF6FC",X"F9FFEF",X"F9FFFD",X"FFFEFF",X"CCD7EB",X"BDCEE0"),
(X"F9FFFF",X"D3FBF0",X"4DDFB0",X"00CC89",X"22D89F",X"36E3AD",X"5DFFD1",X"7CFFDB",X"88FFEC",X"70FED8",X"50E2BD",X"62CDB3",X"E3FFFC",X"FEFAF9",X"F7FEF7",X"F8FFFA",X"FFF7FF",X"F9FCFF",X"CAAAD3",X"833C88",X"550C51",X"4F004D",X"AC4DB5",X"CD87DD",X"F7B5FD",X"FFD0FF",X"FFE1FF",X"E0DCED",X"A3C1B9",X"7EBFA7",X"6BC8AB",X"59C4A8",X"E9F5F5",X"FFFDFF",X"FEFFFF",X"FCFDFF",X"F7F3F2",X"E3FFF6",X"90DBC4",X"256F5E",X"09000A",X"270F25",X"B38EAF",X"FFDBFF",X"FFD5FF",X"FFD9FF",X"FFDBFF",X"FFCDFF",X"9580A7",X"030005",X"342637",X"D0BABD",X"FFF8F2",X"F9FFFD",X"F2F8EA",X"FFF6FF",X"FFFCF3",X"F1FCF8",X"F4FFFF",X"EAEAE2",X"40273A",X"230200",X"794604",X"E39543",X"FFD079",X"FFE18D",X"FFE89D",X"FFDFA3",X"BC9C75",X"100000",X"9A959C",X"FCFDFF",X"FFF6FB",X"EDFFFF",X"92DED4",X"001200",X"070709",X"6D636B",X"F4E5EC",X"FFD5FF",X"FFD0FF",X"FFCEFF",X"DD9CDE",X"770672",X"D5A6EA",X"F1FFFF",X"F5FFF3",X"FFF5FF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FDFDFD",X"FFFCFF",X"F6C3E4",X"1F0000",X"372731",X"1D0F06",X"D8CCC0",X"FEFFE8",X"FFFBFF",X"FFFBF6",X"FFFBFE",X"F8FBFF",X"F9FFFF",X"F9FAFC",X"FEFFFD",X"FBFFFD",X"FBFDFC",X"FFF7FF",X"EEFFFF",X"9DC0D3",X"2C63A3",X"0667B6",X"0F70B7",X"68AEF3",X"A8EEFF",X"C8FFFF",X"C1FAFF",X"ECFCFF",X"ECE9FF",X"A89FB0",X"580E27",X"69081C",X"C9AEA5",X"F8F4F1",X"FBFFFE",X"F1FFFD",X"EAF9F6",X"FFFFFF",X"FFF5FE",X"FFFDFF",X"93A1AC",X"073F94",X"4561AB",X"00060D",X"8C8187",X"E6C7CD",X"FFF4CD",X"FFE4C7",X"BDB5B3",X"676B6E",X"0D0000",X"D2C4C3",X"FFFFFA",X"FFFCFB",X"EFF9F8",X"F4FFFF",X"FFFEFD",X"FDC3D1",X"A30A1E",X"C32323",X"A3000B",X"FFA9C2",X"FEF9FF",X"FEFFFF",X"FFFCF3",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FDFFFE",X"FDFFFE",X"FEFEFE",X"FDFDFD",X"FEFCFD",X"FDFEFF",X"CCCDD1",X"060009",X"B53774",X"BE0053",X"FE93CB",X"FFF8FF",X"FEFFFF",X"FDFCF8",X"FCFAFB",X"FDFDFF",X"F8FAF9",X"FBFDF8",X"FCFEF9",X"FEFFFF",X"BBBAC0",X"000237",X"2992C9",X"4FB9F3",X"B1FBFF",X"DEFCFA",X"F7F1F1",X"CCD2CE",X"ADA5A2",X"0D0004",X"C9C9CB",X"FAFCFF",X"EFEEF6",X"FFFFEF",X"FFFCF3",X"FAFCFF",X"D7F5FF",X"54B1DA",X"3189B1",X"468CAE",X"3C697E",X"84969A",X"ADB2AB",X"D2D8CE",X"D4DFD9",X"B7C0BF",X"ADC5C5",X"8ACCDC",X"39A5CB",X"1882A9",X"AAE3F4",X"F5FFFF",X"FAF6F3",X"F9FFFF",X"FFFFE1",X"F4F180",X"BDD016",X"CEE20F",X"DADE17",X"FEFC81",X"FEFEF2",X"F3FAE8",X"FFFFFA",X"FBFFFF",X"FCFFFF",X"FEF8FF",X"FFFEFF",X"FFF4FD",X"AF6B84",X"620100",X"8D3134",X"58000A",X"EDAABC",X"FCF6F6",X"F3FEFA",X"FFFBFF",X"FFFBFF",X"FFF1FF",X"FC8FC6",X"C20065",X"C40064",X"CC6499",X"FFEBF7",X"FFFDFB",X"FFFEFA",X"F5FBF7",X"FFFDFF",X"FAF4FF",X"FBFFFF",X"F7FCFF",X"F3F5F4",X"EFFFFF",X"93C3C3",X"1A8571",X"008277",X"7AC2B7",X"FFFCF7",X"FCFFFD",X"FEFFFF",X"FFFAFF",X"F1FFF7",X"FFF9FF",X"D8E1E0",X"000405",X"6A5E24",X"D0C52B",X"F1E6A6",X"FFFCF8",X"FFFDFF",X"FFF9FF",X"FFFBFC",X"EFF4EE",X"FFFBFF",X"F5FFFF",X"DAC8D8",X"3F2D3D",X"080007",X"2E002B",X"B86DB0",X"FFBEFF",X"FFCBFF",X"FFCDFF",X"FFD0FF",X"FFC0FF",X"FC94E3",X"DE4EC0",X"9F0774",X"F56ECA",X"FFCEFF",X"FFF5FF",X"F2F7FB",X"FFFCFB",X"FFF3EF",X"FCF6FF",X"FCFFFF",X"FCFFFF",X"FFF2FF",X"B79D9E",X"16000E",X"060013",X"595E5A",X"DBD9DC",X"FFF8FF",X"F2F2FC",X"E9FBFD",X"D5E1F7",X"867EB7",X"090945",X"97B3DA",X"F1FFF8",X"FDFFF2",X"F8F8F0",X"FCFFFF",X"FFFDFF",X"FFF5F5",X"FFFDFF",X"DBF5FF",X"6285E1",X"0850BE",X"004A94",X"628FE4",X"ABC4FF",X"D0F9FF",X"C8F5FF",X"B3DAFF",X"6E82A7",X"BBD5F8"),
(X"F4FDFC",X"BDE5DA",X"23B586",X"00C582",X"11C78E",X"15C28C",X"11B985",X"2CB58B",X"24B388",X"28B690",X"1BAD88",X"5FCAB0",X"E5FFFE",X"FFFEFD",X"F5FCF5",X"F9FFFB",X"FFF6FF",X"F4F7FC",X"FFEEFF",X"FFC4FF",X"CA81C6",X"863184",X"590062",X"510B61",X"54125A",X"521A59",X"36123E",X"01000E",X"000A02",X"105139",X"369376",X"6FDABE",X"F5FFFF",X"FBF6FD",X"FEFFFF",X"FEFFFF",X"FFFCFB",X"EAFFFD",X"BFFFF3",X"93DDCC",X"413342",X"0F000D",X"23001F",X"4A1A44",X"773D70",X"8F528B",X"7B3E79",X"4D114D",X"261138",X"928D94",X"E8DAEB",X"FFF6F9",X"FFFDF7",X"F1FAF5",X"FCFFF4",X"FFF3FF",X"FFFDF4",X"F8FFFF",X"EEF9FD",X"898981",X"14000E",X"74532A",X"B4813F",X"CE802E",X"BA7720",X"CD8C38",X"B98136",X"B28448",X"5E3E17",X"0E0000",X"DDD8DF",X"FAFBFF",X"FFEFF4",X"D9F4EB",X"76C2B8",X"124735",X"000002",X"070005",X"1D0E15",X"4E0D69",X"55165D",X"5C0E4A",X"420143",X"72016D",X"FFD3FF",X"F1FFFF",X"F0FFEE",X"FFF6FF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FDFDFD",X"E5E1F0",X"996687",X"390D0E",X"0A0004",X"100200",X"807468",X"D6DCC0",X"F7F2FF",X"FFFAF5",X"FFFCFF",X"F8FBFF",X"F9FFFF",X"F8F9FB",X"FDFFFC",X"FBFFFD",X"F9FBFA",X"FFF5FF",X"EFFFFF",X"E4FFFF",X"ABE2FF",X"3FA0EF",X"0364AB",X"054B90",X"2A70B6",X"366E91",X"427B98",X"4D5D7F",X"000019",X"04000C",X"994F68",X"FFB7CB",X"FFF1E8",X"FFFEFB",X"F7FBFA",X"F5FFFF",X"F5FFFF",X"FAFAFC",X"FFF7FF",X"F1EEF9",X"5B6974",X"000B60",X"25418B",X"00030A",X"070002",X"3F2026",X"C39D76",X"896E51",X"060000",X"020609",X"655256",X"FDEFEE",X"FEFDF8",X"FCF8F7",X"F8FFFF",X"EDFEF8",X"EEEAE9",X"B87E8C",X"8F000A",X"A60606",X"A5000D",X"AC3A53",X"D7D2D8",X"FCFEFD",X"FFFFF6",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FDFFFE",X"FDFFFE",X"FDFDFD",X"FDFDFD",X"FEFCFD",X"D9DADC",X"3C3D41",X"08000B",X"860845",X"BE0053",X"831850",X"D4C2D2",X"F3F5F4",X"FFFFFB",X"FEFCFD",X"FEFEFF",X"FCFEFD",X"FEFFFB",X"F9FBF6",X"E9EBEA",X"8A898F",X"101D52",X"3099D0",X"1882BC",X"38829D",X"193735",X"040000",X"010703",X"060000",X"1E0A15",X"DFDFE1",X"FCFEFF",X"FFFEFF",X"FFFFEF",X"FFFCF3",X"FAFCFF",X"E8FFFF",X"AEFFFF",X"83DBFF",X"2F7597",X"001126",X"000509",X"000500",X"000400",X"000400",X"000403",X"000707",X"1F6171",X"0F7BA1",X"339DC4",X"C9FFFF",X"F2FFFF",X"FDF9F6",X"F4FDFC",X"F8EDCF",X"D0CD5C",X"C0D319",X"C9DD0A",X"CCD009",X"D1CF54",X"E0E0D4",X"F9FFEE",X"FFFFFA",X"F6FBFE",X"F9FCFF",X"FDF7FF",X"FFFEFF",X"E2CED7",X"56122B",X"600000",X"65090C",X"5D000F",X"A36072",X"ECE6E6",X"F2FDF9",X"FEF4FC",X"FFF9FF",X"E9BFCD",X"8B1E55",X"B9005C",X"C40064",X"760E43",X"A78B97",X"F9F1EF",X"FFFEFA",X"FBFFFD",X"FFFDFF",X"FFFBFF",X"FBFFFF",X"FAFFFF",X"FEFFFF",X"ECFFFF",X"D8FFFF",X"78E3CF",X"007F74",X"7AC2B7",X"FDFAF5",X"F7FCF8",X"FDFFFE",X"FFF4FB",X"F5FFFB",X"FEF4FD",X"6D7675",X"000102",X"493D03",X"AFA40A",X"B8AD6D",X"D7D2CE",X"F3F0F9",X"FFF5FD",X"FFFBFC",X"FCFFFB",X"FFF7FB",X"F7FFFF",X"FFF3FF",X"F2E0F0",X"A597A4",X"A45DA1",X"611659",X"A65598",X"AB599B",X"9F4A8D",X"9B4187",X"B2509B",X"8B2372",X"D646B8",X"D139A6",X"D54EAA",X"DE90CA",X"ECDEF5",X"F5FAFE",X"FFFBFA",X"FFF3EF",X"FFFCFF",X"F1F5F4",X"F8FBFF",X"FFF9FF",X"FFEDEE",X"C0A8B8",X"20132D",X"000200",X"020003",X"524755",X"4E4E58",X"16282A",X"000117",X"010032",X"B0B0EC",X"E4FFFF",X"F2FFF9",X"FAFEEF",X"FFFFF8",X"FCFFFF",X"FCF6FA",X"FFF6F6",X"FBF9FF",X"97B1D2",X"062985",X"0038A6",X"004A94",X"063388",X"0B2474",X"19425E",X"1A4770",X"0E3576",X"00072C",X"C4DEFF"),
(X"FAF8FD",X"DAD9DE",X"C3D6D0",X"C3F3DD",X"C8FEE6",X"CBEFE3",X"C8E1DB",X"C4DFD8",X"BCE0D6",X"BADED4",X"C3E2DA",X"D9EEE9",X"EFF9F8",X"FBFFFF",X"FBFFFF",X"F8FFFF",X"FCF8FF",X"FFFDFF",X"FEF9FF",X"FDF9F8",X"FAF4F4",X"EDDFEC",X"E7CCEB",X"AB87B3",X"8F6398",X"83648E",X"78617E",X"6D556D",X"695E6F",X"ABB4B9",X"D6E0DF",X"F8F4F1",X"FEFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFDFE",X"FFFCFD",X"FCFEFD",X"F5FFFC",X"EAEAF2",X"D4C5D8",X"A481A2",X"8D5E8A",X"90618F",X"7D5780",X"8D708F",X"CDB5CF",X"F5E4FF",X"F9F4FB",X"FAFFF4",X"F9FFFD",X"F8FCFF",X"F9FFF5",X"FAFFF7",X"F8FFFF",X"FEFFFF",X"FFFAFF",X"FFEFF7",X"CFC0C3",X"DDD4CF",X"EBE5D7",X"F0E3D2",X"F3DECB",X"F2D9C3",X"DECCB6",X"E4CEC0",X"E6CBC4",X"D1C3C0",X"D7DCD8",X"F7F8FC",X"FFF8FF",X"FAF9FE",X"DCE8E8",X"C6E1DC",X"D6E1E3",X"EADAE5",X"D8D2DC",X"C9C9D1",X"D7C0D0",X"D5C0D1",X"D5C0D1",X"DCC7D6",X"E7DAE4",X"F6F1F5",X"FEFFFF",X"FEFFFD",X"FFFFFD",X"FEFFFF",X"FEFFFF",X"FEFFFB",X"FFFFFB",X"FFFEFF",X"FFFEFF",X"FEFFFF",X"F8FFFF",X"EEDEE8",X"DACDD6",X"D9CED4",X"E6DDE2",X"DBD5D7",X"C6C0C2",X"D4D0CF",X"F7F6F4",X"FDFCFF",X"FDFDFD",X"FFFCFA",X"FFFEFB",X"F7FFFF",X"FFFFFF",X"FFF9FF",X"F3FFFB",X"FDF9F6",X"F9F9F9",X"F8FDFF",X"F8FFFF",X"F0FBFF",X"CFDDE8",X"9CB3C5",X"7692AA",X"5E88AE",X"6587A3",X"677C8F",X"8E94A4",X"DBD0E0",X"FFF0FF",X"FFF7FF",X"FCFFFF",X"FFFDFA",X"FFFEFF",X"FDFCFF",X"FCFCFE",X"FFFEFD",X"FFFBFA",X"E7E7E9",X"CBCED3",X"CADDE4",X"D3DBE8",X"DED7E7",X"E0D3DA",X"DFD2CA",X"DAD1C0",X"D4CCBF",X"CEC7C1",X"D6C1CA",X"F0DDE3",X"F9FBFA",X"EEFFFF",X"F2FFFF",X"FFF8FF",X"FCF2FB",X"E1EDE9",X"D2C2C5",X"E7CFCF",X"F5D5D6",X"F1CACF",X"E2C1CA",X"E3CFDA",X"F1EEF5",X"F8FFFF",X"FEFFFD",X"FFFEFF",X"FFFCFF",X"FEFEFF",X"FAFFFE",X"FAFFFB",X"FCFDFF",X"F8FDFF",X"E2E2E0",X"D6CACA",X"CAD1C9",X"EBDCDF",X"ECD5DF",X"D0C3CC",X"E7C7D2",X"FAEEEE",X"FFFFFF",X"FFFFFF",X"FCFCFC",X"FAFAFA",X"FFFFFF",X"FCFCFC",X"E6E6E6",X"CCCCCC",X"D3DDE7",X"C9E5E9",X"C1E7EA",X"C0DDE3",X"C5CBD7",X"CBBFCD",X"C9BFC8",X"C6C4C9",X"EBD7E0",X"F9EFF8",X"FBFFFF",X"F4FFFF",X"F4FEFD",X"FCFFFB",X"FFFFFB",X"FDFCFA",X"F7FFFB",X"F3F4F6",X"F0EBF2",X"D4CFD6",X"878586",X"666563",X"635F5E",X"665D60",X"696461",X"5C5F66",X"657283",X"AFBFD6",X"EAF5FF",X"F4F6FF",X"FFFCFF",X"FFF9FE",X"FFFAF1",X"F4E8D8",X"EAE1C4",X"EFE9C7",X"F4F1D2",X"ECECD0",X"DEE0C8",X"D8DAC2",X"F9F8FD",X"FAF9FE",X"FAFBFD",X"FBFCFE",X"FEFEFE",X"F7F5F6",X"E4E0DF",X"D0CACA",X"DFD2DB",X"E9D2DA",X"E1CDCF",X"CDC7C7",X"D7D6DB",X"FCF2FB",X"FFFBFF",X"FBFBFB",X"CDADC5",X"884A6F",X"C16F9D",X"A46487",X"916E82",X"746069",X"E9E0E5",X"FEFEFF",X"FFFFF3",X"FFFFFD",X"FCFFFF",X"FCFFFF",X"FFFEFF",X"FFFDFC",X"FFFCF5",X"FBFDF2",X"E9FFFC",X"C2D7D2",X"B9C5C1",X"F7FDFB",X"FDFFFE",X"FFFFFF",X"F5F7F6",X"FEFFFF",X"EEECEF",X"C8C6C7",X"D7D6D2",X"E5E5DD",X"E7E7DD",X"DBDBD3",X"CCCBC7",X"F1F0EE",X"FAFEFF",X"F3FFFB",X"FFF8F4",X"FFFCF5",X"F8FFFA",X"FBFEFF",X"F4FEFF",X"FFF3FF",X"FAE6EF",X"D6B5D4",X"B281B8",X"A86EAB",X"AD72A8",X"B97EAC",X"C789BA",X"D190C8",X"BF78A4",X"9F5D8B",X"50163C",X"59233D",X"9E678F",X"DAA6E4",X"FCD4FF",X"FFE8FF",X"FFF6FF",X"FFF6FF",X"FFFDFF",X"F9F4F8",X"FFFCFE",X"FFFBFF",X"E1DDEB",X"BABBCD",X"6C6E7A",X"585B64",X"646569",X"615F60",X"B7B3B2",X"EBEAE8",X"F1FAF7",X"F4FFFF",X"F5FFF6",X"FBFFFB",X"FCFFFD",X"FDFCF8",X"FFFEFA",X"FFFFFB",X"E8F1F0",X"C8D7DA",X"D3D8EE",X"D6D8EF",X"CFDAEE",X"C3DAE8",X"BFD3DE",X"C3C9D7",X"C0C7D1",X"B7CACE",X"CFD0D4",X"E7E8EC"),
(X"FFFDFF",X"FDFCFF",X"F2FFFF",X"E0FFFA",X"D7FFF5",X"E3FFFB",X"EDFFFF",X"EAFFFE",X"E7FFFF",X"E4FFFE",X"E5FFFC",X"EFFFFF",X"F8FFFF",X"FBFFFF",X"F6FCFC",X"F3FCFB",X"FEFAFF",X"FCF9FF",X"F9F4FA",X"FFFDFC",X"FFFDFD",X"FFF7FF",X"FFF1FF",X"FFE9FF",X"FFDCFF",X"FFE5FF",X"FFECFF",X"FFF2FF",X"F8EDFE",X"F6FFFF",X"F5FFFE",X"FFFEFB",X"FDFFFE",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FFFDFE",X"FFFCFD",X"FBFDFC",X"F5FFFC",X"F8F8FF",X"FFF8FF",X"FFE9FF",X"FFD9FF",X"FFDEFF",X"FFE3FF",X"FFE8FF",X"FFF2FF",X"FFEFFF",X"FFFBFF",X"FCFFF6",X"FAFFFE",X"FBFFFF",X"FCFFF8",X"FBFFF8",X"F8FFFF",X"FEFFFF",X"FFFCFF",X"FFF7FF",X"FFFAFD",X"FFFDF8",X"FFFFF1",X"FFFBEA",X"FFF5E2",X"FFFAE4",X"FFF5DF",X"FFFAEC",X"FFF8F1",X"FFF3F0",X"F8FDF9",X"FEFFFF",X"FFF9FF",X"FFFEFF",X"F3FFFF",X"E8FFFE",X"F7FFFF",X"FFF9FF",X"FFFBFF",X"FEFEFF",X"FFF6FF",X"FFF2FF",X"FFF0FF",X"FFEFFE",X"FFF6FF",X"FFFDFF",X"FEFFFF",X"FEFFFD",X"FDFCFA",X"FEFFFF",X"FEFFFF",X"FEFFFB",X"FFFFFB",X"FFFEFF",X"FFFEFF",X"FEFFFF",X"F8FFFF",X"FFF4FE",X"FFF9FF",X"FFFBFF",X"FFFCFF",X"FFFCFE",X"FFFCFE",X"FFFDFC",X"FFFEFC",X"FDFCFF",X"FEFEFE",X"FFFCFA",X"FFFEFB",X"F7FFFF",X"FFFFFF",X"FFFAFF",X"F3FFFB",X"FFFDFA",X"FBFBFB",X"F5FAFD",X"F2FCFE",X"F2FDFF",X"EFFDFF",X"E5FCFF",X"DDF9FF",X"D4FEFF",X"E3FFFF",X"E7FCFF",X"F0F6FF",X"FFFAFF",X"FFF7FF",X"FDF2FA",X"F9FDFC",X"FFFDFA",X"FFFEFF",X"FFFEFF",X"FDFDFF",X"FFFDFC",X"FFFEFD",X"FFFFFF",X"F7FAFF",X"EEFFFF",X"F7FFFF",X"FFFBFF",X"FFFAFF",X"FFFCF4",X"FFFEED",X"FFFEF1",X"FFFCF6",X"FFF0F9",X"FFF8FE",X"FEFFFF",X"EFFFFF",X"F1FEFF",X"FFF8FF",X"FFFAFF",X"F5FFFD",X"FFFAFD",X"FFF8F8",X"FFF5F6",X"FFF1F6",X"FFF2FB",X"FFF8FF",X"FFFDFF",X"F7FFFF",X"FEFFFD",X"FFFEFF",X"FFFBFF",X"FEFEFF",X"F9FFFD",X"FAFFFB",X"FBFCFE",X"F8FDFF",X"FCFCFA",X"FFFBFB",X"FBFFFA",X"FFF9FC",X"FFF3FD",X"FFF8FF",X"FFF4FF",X"FFFBFB",X"FDFDFD",X"FFFFFF",X"FDFDFD",X"FBFBFB",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FAFAFA",X"F4FEFF",X"EAFFFF",X"E4FFFF",X"EAFFFF",X"F9FFFF",X"FFF9FF",X"FFFBFF",X"FFFEFF",X"FFEEF7",X"FFF9FF",X"FBFFFF",X"F7FFFF",X"F6FFFF",X"FCFFFB",X"FFFFFB",X"FFFEFC",X"F9FFFD",X"F8F9FB",X"FFFAFF",X"FFFDFF",X"F4F2F3",X"F8F7F5",X"FFFBFA",X"FFF7FA",X"FBF6F3",X"F7FAFF",X"E7F4FF",X"F1FFFF",X"F5FFFF",X"F6F8FF",X"FFFDFF",X"FFF7FC",X"FFFDF4",X"FFFAEA",X"FFFCDF",X"FFFFDF",X"FFFFE3",X"FEFEE2",X"FBFDE5",X"FDFFE7",X"FEFDFF",X"FDFCFF",X"FAFBFD",X"F9FAFC",X"FFFFFF",X"FFFEFF",X"FFFEFD",X"FCF6F6",X"FFFAFF",X"FFF7FF",X"FFF9FB",X"FEF8F8",X"FDFCFF",X"FFFBFF",X"FFFBFF",X"FAFAFA",X"FFE8FF",X"FFDDFF",X"FFD3FF",X"FFD7FA",X"FFE6FA",X"FFEFF8",X"FFF9FE",X"FFFFFF",X"FFFFF3",X"FFFFFD",X"FCFFFF",X"FCFFFF",X"FFFEFF",X"FFFDFC",X"FFFCF5",X"FCFEF3",X"EAFFFD",X"EAFFFA",X"EDF9F5",X"FBFFFF",X"F6F8F7",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FFFEFF",X"FBF9FA",X"FFFFFB",X"FCFCF4",X"FDFDF3",X"FFFFF8",X"FCFBF7",X"FFFFFD",X"FAFEFF",X"F2FFFA",X"FFF7F3",X"FFFBF4",X"F8FFFA",X"FAFDFF",X"F4FEFF",X"FFF3FF",X"FFF8FF",X"FFEAFF",X"FFDBFF",X"FFDAFF",X"FFDAFF",X"FFD8FF",X"FFD7FF",X"FFD8FF",X"FFD7FF",X"FFBFED",X"C98FB5",X"622C46",X"230014",X"562260",X"6E467A",X"CBADC5",X"E6D9E2",X"FFF5FE",X"F5F0F7",X"FFFDFF",X"FFFAFC",X"FFFAFF",X"FFFCFF",X"F1F2FF",X"F2F4FF",X"F6F9FF",X"F3F4F8",X"FAF8F9",X"FFFEFD",X"F9F8F6",X"F9FFFF",X"F0FFFD",X"F8FFF9",X"FBFFFB",X"FCFFFD",X"FDFCF8",X"FFFBF7",X"FFFFFB",X"F7FFFF",X"EDFCFF",X"F8FDFF",X"FBFDFF",X"F5FFFF",X"EDFFFF",X"F0FFFF",X"F8FEFF",X"F8FFFF",X"F1FFFF",X"F9FAFE",X"FEFFFF"),
(X"F2F7FA",X"FDFCFA",X"FFFDFD",X"FEF9FF",X"F7F5FA",X"FEFEFC",X"FBFFFB",X"F2FFFE",X"FCFFFF",X"FAFEFF",X"FAFEFF",X"FEFCFF",X"FFFAFF",X"FFF8FE",X"FFF9FE",X"FFFCFF",X"FBFFFF",X"F7FDF9",X"FBFFF9",X"FFFFFA",X"F4F3EF",X"FFFCFB",X"FAF6F7",X"FCFAFD",X"FDFCF8",X"FFF7F3",X"FCF5ED",X"F8FFF8",X"F2FFFD",X"F4FEFD",X"F4FDFC",X"F0FFFB",X"FFFBFE",X"FBFFFE",X"FAFFFE",X"FFFDFE",X"FFF9FD",X"FFFAFD",X"FDFBFC",X"FDFBFC",X"F5FFFE",X"F6FCFC",X"FBFFFF",X"FBFFFF",X"FAFBFD",X"FFFEFF",X"FFFAFF",X"FFF2FE",X"FFFDFF",X"FFFFF1",X"FDFFED",X"FDFBFE",X"FFF9FF",X"FFFBFF",X"FFFDFA",X"FFFAFA",X"FFFCFB",X"FBFFFD",X"E8F9F3",X"F2FFFD",X"EFF9F1",X"FCF7F1",X"FFFBF4",X"FFF8F1",X"FFFFF4",X"FCFEF1",X"FFFFF6",X"FFFEFA",X"FFFCF9",X"FCFCFA",X"FCFAFB",X"FBF0F6",X"FAF4F6",X"FDFBFC",X"FAFFFE",X"F4FDFC",X"F3F9F9",X"F2FCFB",X"F8FCFF",X"FFF5FF",X"FFFAFF",X"FFF9FF",X"FFF8FF",X"FFF9FF",X"FEFEFF",X"FEFFFF",X"FFFFFD",X"FFFEFD",X"FEFFFB",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFB",X"FFFFF8",X"FFFEFB",X"FFFCFE",X"FFF8FF",X"FFF9FD",X"FFF9FD",X"FEF9FD",X"FEFCFD",X"FFFDFE",X"FBFBFB",X"F6F6F4",X"F7FFFF",X"FFFCFF",X"FCFFFD",X"FCFFFD",X"FFF9FF",X"FFF9FF",X"F8FFFF",X"F5FFFF",X"FBFAF8",X"FBFCFE",X"FAFFFF",X"FAFFFF",X"FAFEFF",X"FAFFFF",X"F8FFFF",X"F4FFFF",X"F8F7FC",X"FBFFFF",X"F7FFFC",X"F2FFFA",X"F3FFFF",X"F5FDFF",X"F7FDFD",X"FBFFFF",X"FFFEFD",X"FFFEFF",X"FFFFFF",X"FEFCFD",X"FCF8F7",X"FCF8F7",X"FAFAFC",X"F8FCFF",X"FAF9FE",X"FFF9FF",X"FCFBFF",X"F4FEFD",X"F5FFF5",X"FFFFF3",X"FFFEF9",X"FDFEFF",X"FCFFFD",X"FFFEFA",X"FAFDF6",X"F3FFF7",X"F7FCF8",X"FFF3F8",X"FFF6F6",X"FDFFF9",X"FAFAFA",X"FBFBF9",X"F9FCF5",X"F6F8F3",X"F6FBF7",X"F9FDFC",X"F8FEFC",X"F6FDF6",X"FDFFFC",X"FEFEFF",X"FEFDFF",X"FEFEFF",X"FEFDFB",X"FFFCF9",X"FDFBFC",X"FBFCFF",X"F5FAFE",X"FFFAFF",X"FEFEFF",X"FFF4FF",X"FFF5FF",X"F7FEFF",X"FBFAFF",X"EAFDF9",X"FBFBFB",X"FDFDFD",X"FDFDFD",X"FAFAFA",X"F9F9F9",X"FAFAFA",X"FCFCFC",X"FDFDFD",X"F9FCFF",X"F5FCFF",X"F6FBFF",X"FCF7FD",X"FFF4F7",X"FFF4F4",X"FCF8ED",X"F4FBEB",X"FCFFFA",X"FAFFFB",X"FCFCFE",X"FFFDFF",X"FFFCFD",X"FFFAFB",X"FFFDFE",X"FEFFFF",X"FBFFFD",X"F9FAFC",X"F9F6FD",X"FFFEFF",X"FCFAFB",X"FFFEFA",X"FFFCFC",X"FFF8FC",X"FEF9F3",X"FEFFFA",X"F5FFF8",X"F3FFF6",X"F5FDF2",X"FDFAF3",X"FFFBFD",X"FFF4FC",X"F3FEFF",X"FAFFFF",X"FEFFFA",X"FFFFF8",X"FCFFF8",X"F9FBF8",X"FEFCFD",X"FFFCFF",X"FEFDFF",X"FFFFFF",X"FDFDFF",X"F8F9FB",X"F9F9F9",X"FCFAFB",X"FFFBFC",X"FDF9F8",X"F6F7F9",X"F9F8F6",X"FAF9F5",X"F9FBF8",X"F9FAFC",X"FBF9FE",X"FBF9FC",X"F9FBFA",X"F4F9FC",X"FEFEFF",X"FBF9FF",X"FBF8FF",X"FFFBFF",X"FFFAFD",X"FFF8FA",X"FEF5F8",X"FFFCFF",X"FFFEFF",X"FEFFFF",X"FEFFFF",X"FFFFFD",X"FFFCFF",X"FEFAFF",X"FCF8FF",X"F9FDFF",X"F8FDFF",X"FAFFFF",X"FCFFFF",X"F7F8FA",X"FFFEFF",X"FFFDFF",X"FFF6FC",X"FDFBFF",X"FBF9FA",X"FEFDF9",X"F8F7F2",X"F8F8F0",X"FEFDF8",X"FAF9F5",X"FAF9F7",X"FFFAFF",X"F5FFFF",X"FFF8FE",X"FAFEFF",X"F7FFFF",X"FFFBFD",X"FCFDF8",X"FFF5F4",X"F8F7FC",X"FFF8FF",X"FFFAFF",X"FFFBFF",X"FFFBF8",X"FEFBF6",X"FFFDFE",X"FFFDFF",X"FFFBFF",X"FCF1FF",X"FFFBFF",X"FCF2F0",X"B1A5A5",X"675764",X"070000",X"090400",X"340829",X"B284A9",X"E9B4E2",X"FFCFFF",X"FFCDFD",X"FFE1FF",X"FFE9FF",X"FFEBFF",X"FFF1FF",X"FFF6FF",X"FFF6FF",X"FFFAFF",X"FFFAFB",X"FFF3F3",X"F7ECEA",X"FFFDFB",X"FFF9FF",X"FFFAFF",X"FEFFFF",X"FCFFFF",X"FDFFFA",X"FDFAF5",X"FFFAFB",X"FFFCFF",X"F1F9FB",X"F6FAFB",X"FAFCF9",X"FAFCF9",X"FDF9FA",X"FFF6FE",X"FEF8FF",X"F8FCFF",X"FEFFFF",X"F8F9FD"),
(X"FBFFFF",X"FCFBF9",X"FFF9F9",X"FFFBFF",X"FFFDFF",X"FFFFFD",X"FBFFFB",X"F2FFFE",X"F8FCFD",X"F8FCFD",X"F8FCFD",X"FCFAFD",X"FFF8FD",X"FFF7FD",X"FFFAFF",X"FFFDFF",X"F8FEFC",X"FBFFFD",X"FAFFF8",X"FAFBF5",X"FCFBF7",X"FFFEFD",X"FFFBFC",X"FDFBFE",X"FFFEFA",X"FFF8F4",X"FFFDF5",X"F6FFF6",X"EEFFF9",X"F8FFFF",X"F9FFFF",X"F4FFFF",X"FFFBFE",X"FCFFFF",X"FBFFFF",X"FFFDFE",X"FFFAFE",X"FFFBFE",X"FEFCFD",X"FEFCFD",X"F8FFFF",X"F0F6F6",X"F3F7F8",X"FCFFFF",X"FAFBFD",X"F8F6FB",X"FFF6FF",X"FFF5FF",X"FFFCFE",X"FDFEEE",X"FBFEEB",X"FCFAFD",X"FFF8FF",X"FFFBFF",X"FFFCF9",X"FFFBFB",X"FFFCFB",X"FBFFFD",X"F4FFFF",X"F2FFFD",X"F5FFF7",X"FDF8F2",X"FFFBF4",X"FFF2EB",X"FDFDF1",X"FBFDF0",X"F8F8EE",X"FBF6F2",X"FDF9F6",X"FCFCFA",X"FDFBFC",X"FFFAFF",X"FFF9FB",X"FFFEFF",X"FBFFFF",X"F6FFFE",X"F8FEFE",X"F8FFFF",X"FBFFFF",X"FFF5FF",X"FDF7FF",X"FEF7FF",X"FFF6FF",X"FEF7FE",X"FBFBFD",X"FBFDFC",X"FEFEFC",X"FFFEFD",X"FEFFFB",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFB",X"FFFFF8",X"FFFEFB",X"FFFCFE",X"FFFCFF",X"FFF9FD",X"FEF8FC",X"FFFDFF",X"FFFEFF",X"F9F7F8",X"FAFAFA",X"FFFFFD",X"F8FFFF",X"FFFCFF",X"FCFFFD",X"FCFFFD",X"FFF9FF",X"FFF9FF",X"F8FFFF",X"F6FFFF",X"FFFFFD",X"FCFDFF",X"F8FDFF",X"F8FDFF",X"F9FDFE",X"F7FCFF",X"F2FBFF",X"EDFAFF",X"FFFEFF",X"FBFFFF",X"F4FFF9",X"EFFEF7",X"EFFEFB",X"F5FDFF",X"FBFFFF",X"FBFFFF",X"FFFDFC",X"FEFCFD",X"FDFDFF",X"FFFEFF",X"FFFEFD",X"FFFCFB",X"FAFAFC",X"F6FAFD",X"FEFDFF",X"FFFBFF",X"FDFCFF",X"F5FFFE",X"F5FFF5",X"FEFEF2",X"FFFDF8",X"FCFDFF",X"F8FDF9",X"F9F8F4",X"F8FBF4",X"F6FFFA",X"FCFFFD",X"FFF7FC",X"FFF6F6",X"FBFEF7",X"FCFCFC",X"FFFFFD",X"FEFFFA",X"FAFCF7",X"F4F9F5",X"F6FAF9",X"FBFFFF",X"FBFFFB",X"FEFFFD",X"FFFFFF",X"FEFDFF",X"FEFEFF",X"FFFEFC",X"FFFDFA",X"FEFCFD",X"FCFDFF",X"FBFFFF",X"FFF8FF",X"FAFAFC",X"FFF8FF",X"FFFAFF",X"F6FDFF",X"FCFBFF",X"F2FFFF",X"FBFBFB",X"FAFAFA",X"FBFBFB",X"FEFEFE",X"FFFFFF",X"FEFEFE",X"FCFCFC",X"FCFCFC",X"FAFDFF",X"F6FDFF",X"F7FCFF",X"FFFAFF",X"FFF8FB",X"FFF8F8",X"FFFCF1",X"F8FFEF",X"FAFFF8",X"F7FCF8",X"FAFAFC",X"FFFDFF",X"FFFCFD",X"FFFBFC",X"FFFCFD",X"FEFFFF",X"F7FDF9",X"FCFDFF",X"FDFAFF",X"FEFCFF",X"FBF9FA",X"F9F8F4",X"FDF7F7",X"FFFBFF",X"FFFAF4",X"FDFFF9",X"F2FDF5",X"F7FFFA",X"FBFFF8",X"FFFFF8",X"FFFBFD",X"FFF0F8",X"F4FFFF",X"F9FFFF",X"FCFFF8",X"FBFCF4",X"FAFDF6",X"FAFCF9",X"FCFAFB",X"FFF6F9",X"F9F8FD",X"FDFDFF",X"FFFFFF",X"FDFEFF",X"FCFCFC",X"FEFCFD",X"FFFBFC",X"FEFAF9",X"FEFFFF",X"FEFDFB",X"FDFCF8",X"FCFEFB",X"FCFDFF",X"FEFCFF",X"FFFEFF",X"FEFFFF",X"FBFFFF",X"F0F0F8",X"FFFDFF",X"FFFDFF",X"FCF6FA",X"FDEEF1",X"FFFBFD",X"FFF7FA",X"FFFCFF",X"FFFEFF",X"FEFFFF",X"FEFFFF",X"FFFFFD",X"FFFCFF",X"FEFAFF",X"FDF9FF",X"FCFFFF",X"F1F6F9",X"F3F9F9",X"FCFFFF",X"FEFFFF",X"FFFEFF",X"FFFDFF",X"FFFBFF",X"FFFEFF",X"FDFBFC",X"FAF9F5",X"FFFFFA",X"FFFFF8",X"FBFAF5",X"FDFCF8",X"FFFFFD",X"FFFAFF",X"F6FFFF",X"FFF9FF",X"FAFEFF",X"F8FFFF",X"FFFBFD",X"FDFEF9",X"FFF6F5",X"FBFAFF",X"FFFAFF",X"FFF9FF",X"FFF9FD",X"FFFAF7",X"FFFCF7",X"FDFBFC",X"FFFAFF",X"FEF3F9",X"FFFAFF",X"FFF6FF",X"FFFAF8",X"FFFBFB",X"F3E3F0",X"B9AEB2",X"6E6956",X"1B0010",X"1C0013",X"8C5785",X"B97BAE",X"A86696",X"C887B1",X"F4BEE2",X"E0B3D4",X"EDD3EE",X"DFC9DE",X"D2C2CF",X"C4B5BC",X"C6B6B7",X"817171",X"9E9391",X"FFFDFB",X"FFF9FF",X"FFF9FF",X"FDFEFF",X"FCFFFF",X"FEFFFB",X"FEFBF6",X"FFF6F7",X"FFF7FA",X"F7FFFF",X"FBFFFF",X"FEFFFD",X"FDFFFC",X"FFFCFD",X"FFF7FF",X"FEF8FF",X"F8FCFF",X"FDFEFF",X"FAFBFF"),
(X"FCFFFF",X"F6FEF3",X"FCFDF8",X"FFFBFF",X"FFF8FF",X"FDF9F6",X"FDFDF5",X"FFFCFF",X"FFFDFF",X"FFFEFF",X"FFFFFF",X"FFFEFF",X"FFFCFF",X"FFFCFF",X"FDFDFF",X"F9FDFE",X"FCFAFB",X"FFFFFD",X"F9F9F7",X"F9F4F8",X"FFFAFF",X"FFF5FF",X"F7F6F2",X"FAFFF3",X"FCFCFF",X"FBF2F7",X"FFFEFB",X"FBFFFA",X"F7FDF9",X"FFF7FA",X"FFF6F7",X"FAF9F5",X"FEFFFF",X"F4FFFF",X"F2FFFF",X"FEFFFF",X"FFFDFF",X"FEFFFF",X"FDFFFE",X"FFFCFE",X"FAFCF9",X"FFFDFE",X"FFFDFF",X"FFFEFF",X"FEFFFF",X"FBFFFD",X"F9FFFD",X"FBFFFD",X"FFFBFF",X"FEFDF8",X"FDFFF4",X"FFFCFF",X"FFFAFF",X"FFFBFF",X"FFFDFF",X"FFFDFF",X"F9FFF8",X"FEFFFA",X"FFF8F9",X"FFF5F9",X"FFFBFF",X"FEFEFF",X"FAFFFE",X"F9FFFF",X"FFFBFF",X"FFFCFF",X"FFFDFF",X"FFFFFF",X"FFFEFF",X"FFFCFF",X"FFFCFD",X"FFFFFD",X"FEFDF9",X"FBFDF8",X"FBFDFA",X"FAFFFB",X"FDFFFC",X"FFFDFC",X"FCFEFD",X"EDFFFC",X"F8FFFF",X"FCFFFF",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FFFEFF",X"FFFCFE",X"FCFFF6",X"FFFFFF",X"FFFCFF",X"FFFDFF",X"FEFFFB",X"FEFFF6",X"FFFDFA",X"FFF8FE",X"F9FAFC",X"FCFDFF",X"FEFFFF",X"FDFEFF",X"FBFDFC",X"FBFDFC",X"FCFEFD",X"FCFEFD",X"FDFEFF",X"FFFCFF",X"F8FFFF",X"F8FFFF",X"FFFDFF",X"FFFEFF",X"FAFFFF",X"FFFAFF",X"FEFFFF",X"FBFFFF",X"F9FDFE",X"FDFDFB",X"FFFFFA",X"FFFEFA",X"FFFEFF",X"FEFFFF",X"FBFBF1",X"FEF9F3",X"FFFBFD",X"FFFAFF",X"FFFAFD",X"FFFEF9",X"FFFFF3",X"FFFFED",X"FFFFFF",X"FEFEFE",X"FCFCFC",X"FFFEFC",X"FFFFFD",X"FFFFFD",X"FFFFFF",X"FEFFFF",X"FEFBF6",X"FFF8F9",X"FDFBFE",X"F5FFFD",X"FBFFFC",X"FFF7FB",X"FFF7FF",X"FFFCFF",X"F1FFFF",X"FDFEFF",X"FFFBFC",X"FFFAF9",X"FFF9F9",X"FFF9FC",X"FFFBFC",X"FBFFFC",X"FBFCFE",X"FBFFFF",X"FAFFFF",X"F8FFFF",X"FAFFFE",X"FEFEFC",X"FFFEF9",X"FFFBF5",X"FFFEFF",X"FCFFFF",X"FBFFFF",X"FFFFFF",X"FFFDFB",X"FFFDFA",X"FFFEFD",X"FEFDFF",X"FFF8FF",X"FFFBFF",X"F9FFFD",X"FCF7FB",X"FFF5FF",X"FFFEFF",X"FFFEFF",X"F0FFFC",X"FFFFFF",X"FDFDFD",X"FBFBFB",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFAFA",X"FFFAFB",X"FFF9FB",X"FFFAFE",X"FFFCFE",X"FDFFFE",X"F9FFFF",X"F7FFFF",X"FAFFF4",X"FEFFF7",X"FFFEFA",X"FFFCFB",X"FFFBFD",X"FFFCFF",X"FFFDFF",X"FAFEFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FDFDFF",X"FFFFFD",X"FEFDF8",X"FFF9F9",X"FFFBFE",X"FAF9FF",X"FDFBFF",X"FDFBFE",X"FFFEFB",X"FFFFF6",X"F8FFF3",X"F5FFFA",X"F2FFFB",X"F8FFFF",X"FCFFFF",X"FEFCFF",X"FEFCFD",X"FCFFFF",X"FCFFFF",X"FFFEFF",X"FFF8FE",X"FEFCFF",X"FEFEFF",X"FFFFFF",X"FEFEFF",X"FEFEFE",X"FFFEFF",X"FFFEFF",X"FFFEFF",X"FFFAFE",X"FFFEFD",X"FFFFFD",X"FFFEFF",X"FFFDFE",X"FDFDFD",X"F8FCFB",X"F6FAF9",X"FFFFFA",X"FEFFFD",X"FFFFFF",X"FFFEFF",X"FDFDFB",X"F9FFFB",X"F2FFF8",X"F1FFF9",X"FFFCFF",X"FFFEFF",X"FFFFFF",X"FFFFFA",X"FFFFFA",X"FFFEFC",X"FFFCFF",X"FDFBFF",X"F9FEFF",X"FBFFFF",X"FCFFFF",X"FBFFFF",X"FAFEFF",X"FEFFFF",X"FEFFFF",X"FEFFFF",X"FCFAFF",X"FFFEFF",X"FEFDFB",X"FDFCF8",X"FDFCF8",X"FEFDFB",X"FFFEFF",X"FCFAFB",X"FFF8FE",X"FFFDFF",X"FEFDFF",X"F7FFFF",X"FEFDFF",X"FFF9FE",X"FAFFF7",X"FAFFF2",X"FDFCF8",X"FFFEF9",X"FFFFF5",X"FDFFF4",X"FDFFF9",X"FCFFFD",X"FAFFFF",X"F4FCFE",X"F8FFF8",X"F4FEFF",X"F5FEFF",X"F8FFFE",X"FBFFFD",X"FCFFFF",X"FCFFFB",X"EEF5E3",X"D7DFD2",X"8E888C",X"72516E",X"924F85",X"882B72",X"B64998",X"7F105C",X"841A62",X"8D1251",X"94416F",X"17000F",X"0D1D1A",X"456556",X"B6CDBD",X"EFEFE7",X"FFF8F3",X"FFFAFF",X"FFFCFF",X"FCFDFF",X"F9FEFF",X"FAFFFF",X"FFFFFF",X"FFFDFF",X"FFFAFF",X"FDFDFB",X"FDFFFC",X"FDFFFE",X"FFFEFF",X"FFFDFF",X"FBFFFF",X"F9FFFF",X"F9FFFF",X"FAF9FE",X"FCFBFF"),
(X"FCFFFF",X"FBFFF8",X"FFFFFB",X"FFFBFF",X"FFF9FF",X"FFFEFB",X"FFFFF8",X"FFFDFF",X"FFFAFE",X"FEFCFF",X"FDFDFF",X"FEFCFF",X"FFFCFF",X"FFFDFF",X"FFFFFF",X"FAFEFF",X"FFFEFF",X"FAFAF8",X"FFFFFD",X"FEF9FD",X"FFF4FE",X"FFF4FE",X"FFFFFB",X"F3FBEC",X"FCFCFF",X"FFF8FD",X"FCF7F4",X"FBFFFA",X"FBFFFD",X"FFFCFF",X"FFFBFC",X"FFFFFB",X"FEFFFF",X"F4FFFF",X"F2FFFF",X"FEFFFF",X"FFFDFF",X"FEFFFF",X"FEFFFF",X"FFFDFF",X"FEFFFD",X"FFFEFF",X"FFFDFF",X"FCF8F9",X"FBFDFC",X"F8FEFA",X"F5FEF9",X"FBFFFD",X"FFFCFF",X"FFFEF9",X"FFFFF6",X"FFFDFF",X"FFFAFF",X"FFF9FF",X"FFFAFF",X"FDFBFF",X"F7FEF6",X"FAFBF6",X"FFF7F8",X"FFFBFF",X"FFFCFF",X"FFFFFF",X"F6FCFA",X"F9FFFF",X"FEF7FF",X"FFFBFF",X"FFFDFF",X"FEFEFF",X"FFFEFF",X"FFF9FC",X"FFF7F8",X"FEFDFB",X"FFFFFB",X"FEFFFB",X"FEFFFD",X"FCFFFD",X"FDFFFC",X"FCF8F7",X"F9FBFA",X"F0FFFF",X"F6FFFF",X"F9FDFE",X"FCFCFE",X"FEFEFF",X"FEFFFF",X"FEFFFF",X"FFFEFF",X"FFFDFF",X"FCFFF6",X"FFFFFF",X"FFFCFF",X"FFFDFF",X"FEFFFB",X"FEFFF6",X"FFFDFA",X"FFF8FE",X"FCFDFF",X"FEFFFF",X"FEFFFF",X"FBFCFE",X"FDFFFE",X"FEFFFF",X"FEFFFF",X"FCFEFD",X"FDFEFF",X"FFFDFF",X"F8FFFF",X"F8FFFF",X"FFFDFF",X"FFFEFF",X"FBFFFF",X"FFFAFF",X"FAFBFD",X"FBFFFF",X"FCFFFF",X"FFFFFD",X"FFFFFA",X"FFFBF7",X"FDFBFC",X"FBFCFF",X"FEFEF4",X"FFFCF6",X"FFFBFD",X"FFFAFF",X"FFFBFE",X"FEFDF8",X"FFFFF2",X"FFFCE9",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFD",X"FDFCFA",X"FAF9F7",X"FAFAFA",X"FBFCFE",X"FFFFFA",X"FFFBFC",X"FFFEFF",X"F7FFFF",X"FCFFFD",X"FFF9FD",X"FFF8FF",X"FFFDFF",X"F0FFFF",X"FEFFFF",X"FFFCFD",X"FFF8F7",X"FFF6F6",X"FFF8FB",X"FFFCFD",X"FAFFFB",X"FBFCFE",X"F9FDFE",X"F9FFFF",X"F9FFFF",X"FBFFFF",X"FFFFFD",X"FFFFFA",X"FFFEF8",X"FFFEFF",X"FCFFFF",X"FBFFFF",X"FFFFFF",X"FFFDFB",X"FFFDFA",X"FFFEFD",X"FFFEFF",X"FFF9FF",X"FFFBFF",X"FBFFFF",X"FFFCFF",X"FFF8FF",X"FFFEFF",X"FFFEFF",X"EFFFFB",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FBFBFB",X"F9F9F9",X"FAFAFA",X"FDFDFD",X"FFFDFD",X"FFFCFD",X"FFFBFD",X"FFFAFE",X"FFFAFC",X"FAFCFB",X"F5FEFB",X"F4FFFE",X"FAFFF4",X"FFFFF8",X"FFFEFA",X"FFFAF9",X"FFF8FA",X"FFFCFF",X"FFFEFF",X"FCFFFF",X"FCFCFC",X"FCFCFE",X"FDFCFF",X"F9F9FB",X"FFFFFD",X"FEFDF8",X"FFFCFC",X"FFFCFF",X"FEFDFF",X"FFFDFF",X"FFFEFF",X"FFFCF9",X"FBFBF1",X"F8FFF3",X"F4FFF9",X"F1FFFA",X"F6FFFF",X"FBFFFF",X"FFFDFF",X"FFFDFE",X"FBFFFF",X"FCFFFF",X"FFFEFF",X"FFF9FF",X"FFFEFF",X"FFFFFF",X"FEFEFF",X"FEFEFF",X"FEFEFE",X"FEFCFD",X"FDFBFC",X"FDF9FA",X"FFF7FB",X"FFFDFC",X"FFFFFD",X"FFFCFD",X"FFFEFF",X"FFFFFF",X"FCFFFF",X"FBFFFE",X"FCFBF6",X"FEFFFD",X"F7F7F9",X"FEFCFF",X"FAFAF8",X"F9FFFB",X"F2FFF8",X"F5FFFD",X"FFFCFF",X"FFFEFF",X"FFFFFF",X"FFFFFA",X"FFFFFA",X"FFFFFD",X"FFFCFF",X"FEFCFF",X"F8FDFF",X"FBFFFF",X"FCFFFF",X"F9FDFF",X"F7FBFE",X"FBFCFF",X"FDFEFF",X"FCFDFF",X"FFFDFF",X"FFFEFF",X"FFFFFD",X"FEFDF9",X"FDFCF8",X"FFFFFD",X"FFFEFF",X"FCFAFB",X"FFF8FE",X"FFFDFF",X"FFFEFF",X"F8FFFF",X"FEFDFF",X"FFF9FE",X"FBFFF8",X"FBFFF3",X"FFFFFB",X"FFFFFA",X"FFFFF6",X"FCFEF3",X"FBFEF7",X"FBFFFC",X"FBFFFF",X"F9FFFF",X"F8FFF8",X"F8FFFF",X"F8FFFF",X"F9FFFF",X"F2F8F4",X"FCFFFF",X"FAFFF9",X"FCFFF1",X"FBFFF6",X"FDF7FB",X"FFE0FD",X"F3B0E6",X"FDA0E7",X"FFA8F7",X"FF98E4",X"FE94DC",X"FF93D2",X"FEABD9",X"DBC0D3",X"E0F0ED",X"EAFFFB",X"F1FFF8",X"FFFFF8",X"FFF8F3",X"FFF7FF",X"FFFCFF",X"FEFFFF",X"FAFFFF",X"F9FFFF",X"FFFFFF",X"FFFDFF",X"FFFAFF",X"FCFCFA",X"FBFDFA",X"FCFEFD",X"FEFCFD",X"FFFDFF",X"FBFFFF",X"F9FFFF",X"F9FFFF",X"FFFEFF",X"FFFEFF"),
(X"FDFDFB",X"F7FDF9",X"F7FDFB",X"FCFAFF",X"FCFAFF",X"FEFFFF",X"FFFFFD",X"FEF8FA",X"FEFFFF",X"FBFFFF",X"F9FFFF",X"FBFFFF",X"FDFEFF",X"FFFFFF",X"FBFFFF",X"F6FFFE",X"FFFBFF",X"F4F4F2",X"FCFFFB",X"FDFFFE",X"FDF5FF",X"FFFAFF",X"EFE9ED",X"BCBBB6",X"C89DCA",X"FFF4FF",X"FFF8FF",X"FFF9FF",X"FFFBFF",X"FBFFFF",X"F4FFF9",X"FBFCF6",X"FFFDFF",X"FFFDFF",X"FFFDFF",X"FFFEFF",X"FBFFFF",X"F8FFFF",X"FBFFFF",X"FFFEFF",X"FDFDF5",X"FFFAF8",X"FFF7FE",X"FFF9FF",X"FFFBFF",X"FCFBFF",X"F8FDF9",X"FBFFFA",X"FFFBFF",X"FDFCFF",X"FCFDFF",X"FDFDFF",X"FEFDFF",X"F8FCFB",X"F3FEF6",X"F0FFF6",X"FBF9FA",X"FFFFFF",X"FCFFFF",X"E1E9EB",X"B6C2C2",X"CCD8D8",X"F8FFFF",X"F8FFFF",X"FCFFFF",X"FEFEFF",X"FCFFFF",X"F8FFFF",X"FBFFFF",X"FFFEFF",X"FFFFFF",X"F9FFFF",X"FCFBF9",X"FFF8F9",X"FFFAFB",X"FAFFFE",X"F3FFFD",X"FFF9FC",X"FFF7FF",X"FFFCFF",X"F8FFFD",X"FCFFFD",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FCFFFF",X"FEFEFE",X"FEFCFD",X"FCFFFA",X"FFFEFF",X"FFFCFF",X"FEFEFF",X"F9FFFF",X"F9FFFF",X"FFFFFF",X"FFFAFF",X"FCFFFF",X"FAFEFF",X"F9FAFC",X"FBFCFE",X"FDFDFD",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"F8FFFF",X"FFFEFF",X"FFFCFF",X"F7FFFD",X"F5FFFD",X"FFFEFF",X"FFFBFF",X"FFFFFF",X"FEFFFF",X"FEFFFF",X"FDFDFB",X"FFFAF6",X"FFFAF7",X"FFFEFF",X"FFFEFF",X"F4FFFF",X"F7FEFF",X"FCF9FF",X"FFF6F9",X"FFFDF9",X"F8FFFD",X"F9FFFF",X"FFFBFF",X"F6FBFF",X"FCFDFF",X"FFFFFD",X"FFFEFB",X"FFFFFD",X"FFFFFF",X"FFFFFF",X"FFFFFD",X"FBFFFB",X"FFFBFC",X"FFFBFE",X"FBFFFF",X"FFFEFF",X"FFF5FE",X"FFF7FF",X"F1FFFF",X"FEFBFF",X"FFFBFF",X"FFFDFF",X"F9FFFF",X"F5FFFF",X"F8FFFF",X"FEFFFF",X"FFFCFF",X"FEFFFF",X"FFFEFF",X"FFFBFF",X"FFF8FF",X"FFF5FE",X"FFF5FB",X"FFF9FB",X"FFFDFE",X"FFFCFF",X"FBFFFF",X"F7FFFF",X"FFFFFD",X"FFFEFA",X"FFFFFA",X"FEFFFD",X"FFFFFF",X"FFFFFD",X"FDFCF7",X"F9FEF7",X"FEFFFA",X"FEFFFD",X"FBFDFA",X"FFF9F6",X"FFFEF4",X"FAFAFA",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFAFB",X"FFFAFA",X"FFFCF9",X"FBFFFA",X"F6FFFA",X"F8FFFF",X"FFFEFF",X"FFFAFF",X"FFF8FE",X"FFFAFD",X"FFFCF9",X"FBFDF8",X"F9FFFB",X"F9FFFF",X"FBFFFF",X"FEFFFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"FCFEFD",X"FFFFFB",X"FCFBF6",X"FFFFFD",X"FFFDFF",X"F7FFFF",X"FCFDFF",X"FFFCFF",X"FFF9FF",X"FFFCFF",X"FFFDFF",X"FFFFFF",X"FDFEF9",X"FFFFFB",X"FFFDFD",X"FFFCFF",X"FFFDFF",X"FEFFFF",X"F7FFFB",X"F7FFFB",X"FAFFFE",X"FDFBFE",X"FDFBFE",X"FDFDFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FFFFFF",X"FBFFFF",X"FBFFFF",X"FDFBFE",X"FFFBFC",X"FDFFFC",X"FCFFFF",X"FFFEFF",X"FBFFF8",X"F2FFF6",X"F8FFFF",X"FFFEFF",X"FFFCFD",X"FBF5F5",X"FFFAFD",X"FFFAFF",X"FCFFFA",X"FEFFF8",X"FFFFFA",X"FFFEFB",X"FFFFFD",X"FFFFFD",X"FFFFFB",X"FFFFF8",X"FCFFFF",X"FDFFFE",X"FEF9FD",X"FFFDFF",X"FFFDFF",X"FFFEFF",X"F9FFFF",X"F8FFFF",X"FFFEFF",X"FEFCFF",X"FFFDFE",X"FFFFFD",X"FFFEFC",X"FCFAFB",X"FBF9FC",X"FFFEFF",X"EBFFF1",X"FFFFF5",X"FFFBFB",X"FEFFFF",X"FDFFFE",X"FDFEFF",X"F8FFFF",X"FEFFFF",X"FCFBF7",X"FEFDF9",X"FFFEFF",X"FFFDFF",X"FFFAFF",X"FFF8FF",X"FFF8FE",X"FFF9F7",X"FFFBF0",X"FFFCFD",X"FFF4FF",X"FFFAFF",X"FEF9FF",X"FCF9FF",X"FEFCFF",X"FCFAFF",X"FBFCFE",X"FCFDFF",X"FFFEFF",X"FFF8FF",X"F9ECFF",X"FFF7FF",X"FEFEFF",X"F4FEFF",X"F8FCFF",X"F4F8FF",X"FFFEFF",X"FFFCFF",X"FFF2F5",X"FFF5F6",X"FFFBF9",X"FFFDF8",X"F1FFF4",X"F8FFF8",X"FCFFFB",X"FEFFFF",X"FEFFFF",X"FBFEFF",X"FAFEFF",X"F9FDFE",X"FFFEF8",X"FFFFFB",X"FFFEFF",X"FFFDFF",X"FFFDFC",X"FEFFF7",X"FFFFF0",X"FFFCEB",X"FFFEFC",X"FEFDFB"),
(X"FFFFFD",X"F8FEFA",X"FBFFFF",X"FFFEFF",X"FFFDFF",X"FBFDFC",X"FFFFFD",X"FFFDFF",X"FAFBFD",X"FAFFFF",X"F9FFFF",X"F8FEFE",X"FAFBFD",X"FDFDFF",X"FCFFFF",X"F9FFFF",X"FEF7FE",X"FFFFFD",X"F6FBF5",X"F8FAF9",X"FFFBFF",X"CEC2CE",X"393337",X"010000",X"3E1340",X"F6DDFB",X"FFFAFF",X"FFF5FC",X"FFF6FA",X"FAFFFE",X"F8FFFD",X"FEFFF9",X"FFFDFF",X"FFFDFF",X"FFFDFF",X"FFFEFF",X"FBFFFF",X"F8FFFF",X"FBFFFF",X"FFFEFF",X"FFFFF8",X"FFFBF9",X"FFFAFF",X"FFF9FF",X"FFF7FF",X"FFFEFF",X"FCFFFD",X"F7FEF6",X"FFFCFF",X"FCFBFF",X"FAFBFF",X"FCFCFF",X"FEFDFF",X"FAFEFD",X"F5FFF8",X"F2FFF8",X"FFFDFE",X"FBFBFD",X"B9BDBE",X"363E40",X"000404",X"475353",X"ECF6F7",X"F9FFFF",X"FCFFFF",X"FBFBFF",X"FBFEFF",X"F8FFFF",X"FAFFFF",X"FFFEFF",X"FFFFFF",X"F7FFFD",X"FFFFFD",X"FFFCFD",X"FFFBFC",X"F8FEFC",X"F4FFFE",X"FFFCFF",X"FFF7FF",X"FFF9FC",X"F7FFFC",X"FBFFFC",X"FEFEFE",X"FEFEFE",X"FDFFFE",X"FBFFFE",X"FFFFFF",X"FFFEFF",X"FCFFFA",X"FFFEFF",X"FFFCFF",X"FEFEFF",X"F9FFFF",X"F9FFFF",X"FFFFFF",X"FFFAFF",X"F6FAFB",X"FCFFFF",X"FEFFFF",X"FEFFFF",X"FCFCFC",X"FEFEFE",X"FFFFFF",X"FEFEFE",X"FFFEFF",X"F8FFFF",X"FFFEFF",X"FFFCFF",X"F7FFFD",X"F5FFFD",X"FFFEFF",X"FFFBFF",X"FFFFFF",X"FDFEFF",X"FDFEFF",X"FFFFFD",X"FFFEFA",X"FFFDFA",X"FFFCFD",X"FAF9FE",X"F1FEFF",X"F8FFFF",X"FFFDFF",X"FFF9FC",X"FFFDF9",X"F6FFFB",X"F7FEFF",X"FFFBFF",X"FBFFFF",X"FEFFFF",X"FEFDFB",X"FFFBF8",X"FFFEFC",X"FFFFFF",X"FFFFFF",X"FBFBF9",X"FBFFFB",X"FFFAFB",X"FFFAFD",X"FBFFFF",X"FFFEFF",X"FFF6FF",X"FFFAFF",X"F4FFFF",X"FFFDFF",X"FFF9FF",X"FDFAFF",X"F8FFFF",X"F5FFFF",X"F7FFFF",X"FBFCFF",X"FCF9FF",X"FEFFFF",X"FEFCFF",X"FFF8FF",X"FFF9FF",X"FFFAFF",X"FFFBFF",X"FFFDFF",X"FFFDFE",X"FFFCFF",X"FBFFFF",X"F7FFFF",X"FFFFFD",X"FFFEFA",X"FFFFFA",X"FEFFFD",X"FFFFFF",X"FFFFFD",X"FEFDF8",X"F9FEF7",X"FCFFF8",X"FEFFFD",X"FEFFFD",X"FFFDFA",X"FFFEF4",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FCFCFC",X"FDFDFD",X"FFFFFF",X"FFFFFF",X"FCFCFC",X"FFFEFF",X"FFFCFC",X"FFFDFA",X"FBFFFA",X"F6FFFA",X"F7FFFE",X"FEFDFF",X"FFF8FF",X"FFFBFF",X"FFFBFE",X"FFFDFA",X"FEFFFB",X"FBFFFD",X"F9FFFF",X"FAFFFF",X"FCFEFD",X"FFFEFF",X"FBFBFD",X"FDFEFF",X"F9FBFA",X"FFFFFB",X"FFFFFA",X"FFFFFD",X"FCFAFF",X"F9FFFF",X"FBFCFF",X"FFFDFF",X"FFFBFF",X"FFFBFF",X"FCF9FF",X"FAFAFC",X"FFFFFB",X"FFFFFB",X"FFFAFA",X"FFF9FE",X"FFFDFF",X"FEFFFF",X"F9FFFD",X"F9FFFD",X"FBFFFF",X"FFFEFF",X"FFFDFF",X"FCFCFE",X"FBFBFD",X"FBFBFB",X"FCFCFC",X"FEFCFD",X"FFFEFF",X"FDFDFD",X"F9FFFF",X"FBFFFF",X"FFFEFF",X"FFFEFF",X"FDFFFC",X"FCFFFF",X"FFFEFF",X"F9FFF6",X"F7FFFB",X"F5FFFC",X"FAF8FB",X"FFFCFD",X"FFFDFD",X"FFFAFD",X"FFF9FF",X"FCFFFA",X"FEFFF8",X"FFFFFA",X"FFFEFB",X"FFFFFD",X"FFFFFD",X"FFFFFB",X"FFFFF8",X"F6FAF9",X"FEFFFF",X"FFFCFF",X"FFFDFF",X"FFFDFF",X"FFFEFF",X"F8FEFE",X"F8FFFF",X"FEFCFF",X"FDFBFE",X"FFFEFF",X"FEFDFB",X"FEFDFB",X"FFFEFF",X"FEFCFF",X"FFFEFF",X"EBFFF1",X"FFFFF5",X"FFFAFA",X"FDFFFE",X"FCFEFD",X"FCFDFF",X"F8FFFF",X"FEFFFF",X"FFFFFB",X"FDFCF8",X"FBF9FA",X"FFFAFF",X"FFF9FF",X"FFF8FF",X"FFFAFF",X"FFFCFA",X"FFFDF2",X"FFF8F9",X"FFF9FF",X"FFF4FF",X"FFFDFF",X"FFFDFF",X"FEFCFF",X"FEFCFF",X"F9FAFC",X"FCFDFF",X"FCFBFF",X"FFF8FF",X"FFF8FF",X"FFF9FF",X"F4F4FC",X"F8FFFF",X"F6FAFF",X"FBFFFF",X"F2F1F7",X"FFFBFF",X"FFF9FC",X"FFF7F8",X"FFFCFA",X"FEFBF6",X"F5FFF8",X"F7FFF7",X"F9FEF8",X"FCFEFD",X"FEFFFF",X"FCFFFF",X"FBFFFF",X"FBFFFF",X"FFFEF8",X"FFFFFB",X"FFFDFE",X"FFFCFE",X"FFFDFC",X"FEFFF7",X"FFFFF0",X"FFFCEB",X"FEFDFB",X"FFFEFC"),
(X"FFFEFA",X"FFFCFF",X"FFFAFF",X"FFF9FF",X"FFF6FE",X"FFFBFF",X"FEFEFF",X"F7FDFB",X"F5F9FA",X"FBFFFF",X"F8FFFF",X"F7FBFC",X"FFFDFF",X"FFF6FB",X"FFFCFF",X"FFFBFF",X"FFF7FF",X"FFFCFF",X"FFFDFF",X"F2F1F6",X"8E8B92",X"07000A",X"514053",X"9F879F",X"D9C9E4",X"F2F6FF",X"F3FFFB",X"FDFEF9",X"FFFEFB",X"FDFDFD",X"F9F9FB",X"FFFCFF",X"FAFFFF",X"FFFCFF",X"FFFBFF",X"F1F5F6",X"F7FFFF",X"FFFFFF",X"FFF6FD",X"FFF8FF",X"FFFAFF",X"FFFBFF",X"FEFDFF",X"F6FEFF",X"F7FFFF",X"FBFFFF",X"FFF9FD",X"FFF8FF",X"FCFEF0",X"FEFFFB",X"FEFFFF",X"FFFDFF",X"FFFAFF",X"FFFBFF",X"FFF6F7",X"FFFDF7",X"F9EDFB",X"9B909E",X"554D58",X"746A73",X"B6ABB3",X"E1D6DC",X"FEF8FC",X"FFFEFF",X"FFFCFF",X"FFF7FB",X"FFFAFF",X"FFFBFF",X"FBF9FC",X"FAFFFF",X"F9FFFF",X"F8FFFF",X"F0FFFF",X"F2FCFD",X"F7FFFF",X"F1FFFF",X"F8FFFF",X"FFFAFF",X"FFFBFF",X"F3FFFF",X"FDFFFC",X"FFFEFD",X"FFFDFD",X"FFFBFB",X"FEFEFE",X"FCFFFF",X"FCFFFF",X"FEFFFF",X"FEFFFF",X"FBFBFB",X"FFFFFD",X"FFFFFD",X"F5F5F7",X"FCFFFF",X"F9FEFF",X"F7FEFF",X"FEFFFF",X"FDFDFD",X"FEFEFE",X"FFFEFF",X"FEFCFF",X"FEF9FD",X"FFFCFF",X"FFFDFF",X"FFF6F7",X"FFFFFF",X"FFF9FF",X"FFF6FC",X"FCFFF6",X"FEFFF6",X"FFFFFA",X"F7FFFF",X"FFFEFB",X"FFFEFF",X"FEFFFF",X"FFFFFF",X"FBFAF8",X"F9F9FB",X"FBFFFF",X"F5FDFF",X"FFFDF1",X"FFFFF8",X"FAFEFD",X"FEFEFF",X"F7FFFD",X"EEFFFF",X"F6FFFF",X"FFF6FF",X"F5FFFF",X"F9FEFF",X"FFFFFB",X"FFFCF9",X"FFFFFF",X"FEFFFF",X"F9F9F9",X"FFFEFA",X"FAFBFF",X"FFFBFF",X"FFFDFF",X"F6FFFF",X"F6FFFF",X"FFFEFF",X"FCF8F5",X"FAFFF7",X"FFFDFA",X"FFFDFE",X"FFFBFF",X"FFF9FF",X"FFFEFB",X"F8FBF4",X"FAFEFD",X"FCFDFF",X"FFFCFA",X"FFFAFE",X"FFFCFF",X"FFFDFF",X"F8F8FA",X"FEFFFF",X"FCFFFF",X"F9FDFF",X"FFFAFF",X"F8FEFE",X"F8FFFF",X"FFFFFD",X"FEFFF9",X"F2FFF5",X"FBFFFF",X"FFFAFF",X"F4FFFF",X"FCFAFD",X"FFF8FF",X"FFF8FF",X"FEFFFF",X"F7FFFF",X"F9FFFD",X"FEFBF4",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FEFEFE",X"FDFDFD",X"F8FFFF",X"FCFFFF",X"FEFFFD",X"F9FFFA",X"EDFFF3",X"F4FFFF",X"F8FFFF",X"FFFEFF",X"F3FEFF",X"F9FFFF",X"FBFFFF",X"F8FCFB",X"F9FFFF",X"F8FFFF",X"F6FAF9",X"FFFFFB",X"FFFDFF",X"FEFEFF",X"FBFFFF",X"FEFFFD",X"F9F8F3",X"FFFFFB",X"FCFFFF",X"F7FFFF",X"FFFCF4",X"FFFCF3",X"FFF7EC",X"FFFFF8",X"FEFFFF",X"FDFDFF",X"FFF7FF",X"FFF9FF",X"FEFFFF",X"F9FAFF",X"FFFBFF",X"FFFAFF",X"FFF9FF",X"FFF2F7",X"FFFDFF",X"FAFDFF",X"FFFEFF",X"FCFAFB",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FDFBFE",X"F7FFFF",X"FEFEFF",X"FFF6FF",X"FFF7FF",X"FFFFFF",X"F9FEF8",X"FEFDFB",X"FFFAFF",X"FCFBF7",X"FFFDFF",X"FEF4FD",X"FFFCFF",X"F9F7FC",X"FFFDFF",X"FFF9FF",X"FFF6FF",X"EFFEF9",X"FBFFFB",X"FFFFF8",X"FFFEFB",X"FFFEFF",X"FCFCFF",X"FFFEFF",X"FEFCFF",X"FFF8F8",X"FFFBFB",X"FCF6F6",X"FFFEFF",X"FBFBFB",X"FBF9FA",X"FFFDFF",X"FFFBFC",X"FEFEFF",X"FEFEFF",X"FEFEFF",X"FEFEFF",X"FEFEFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"F2FFFF",X"FFF8FE",X"F4FDFC",X"F1FFFD",X"FFFDF7",X"FFF5F5",X"FFFCFF",X"FDFCFF",X"FCFFFF",X"FAFFFF",X"F8FFFF",X"FBFFFF",X"FFFEFF",X"FFFEFF",X"F9FFFF",X"F2FFFC",X"FBFFFF",X"FDFBFF",X"FFF6FD",X"FFFAFF",X"FFFCFF",X"FAF6F5",X"FFFEFF",X"FFFAFF",X"FFF6FF",X"FFFDFF",X"F4FAF6",X"FBFFF5",X"FDFDF5",X"FAF5F2",X"FFFBF9",X"FFFDFA",X"FFFFFF",X"F8FCFD",X"F7FFFD",X"F4FDFA",X"FCFFFF",X"F4F5F7",X"FBFFFF",X"F5FDFF",X"F5FFFD",X"F1F8F0",X"FFFFFA",X"FFFFFD",X"FCFCFE",X"FEFEFC",X"FEFAEF",X"FFFFEC",X"F0FFFB",X"F7FFFB",X"FFFFFB",X"FEF8F8",X"FEFCFD",X"FCFFFF",X"FBFBFF",X"FEFCFF",X"F8F8F0",X"FFFFF8"),
(X"FFFFFB",X"FFFBFF",X"FFF4FF",X"FFFBFF",X"FFFBFF",X"FCF6FF",X"FEFEFF",X"FBFFFF",X"FCFFFF",X"F0F6F6",X"F9FFFF",X"F9FDFE",X"FBF6FA",X"FFFAFF",X"FFF9FE",X"FFFDFF",X"FFF9FF",X"FFFCFF",X"FDFBFF",X"F5F4F9",X"B0ADB4",X"D3C8D6",X"FFF1FF",X"FFF4FF",X"FFF7FF",X"FBFFFF",X"F7FFFF",X"FFFFFB",X"FFFBF8",X"FFFFFF",X"FFFFFF",X"FFF8FB",X"F8FEFE",X"FFF7FC",X"FFFBFF",X"FCFFFF",X"F6FFFF",X"FBFBFD",X"FFFAFF",X"FFF9FF",X"FFF5FF",X"FFFAFF",X"F6F5FA",X"F9FFFF",X"F7FFFF",X"F4FAFA",X"FFFBFF",X"FFF6FF",X"FBFDEF",X"F9FBF6",X"FCFDFF",X"FFFDFF",X"FFF7FF",X"FFF8FF",X"FFFCFD",X"FFFCF6",X"F7EBF9",X"D5CAD8",X"FFFBFF",X"FFF8FF",X"FFF8FF",X"FFF5FB",X"FFFDFF",X"FEFCFD",X"FFF6F9",X"FFFBFF",X"FFF5FC",X"FFF7FD",X"FFFEFF",X"F1F6F9",X"F9FFFF",X"F3FDFE",X"F4FFFF",X"F8FFFF",X"F7FFFF",X"EEFFFF",X"F3FBFD",X"FFF4FD",X"FFF9FF",X"F4FFFF",X"FCFEFB",X"FFFCFB",X"FFFCFC",X"FFFCFC",X"FFFFFF",X"FCFFFF",X"FCFFFF",X"FDFFFE",X"FEFFFF",X"FEFEFE",X"FDFCFA",X"F8F7F5",X"FFFFFF",X"FCFFFF",X"F9FEFF",X"F9FFFF",X"FEFFFF",X"FBFBFB",X"FDFDFD",X"FFFEFF",X"FFFEFF",X"FFFDFF",X"FFFDFF",X"FFFBFF",X"FFFCFD",X"FFFFFF",X"FFF9FF",X"FFF9FF",X"FEFFF8",X"FDFFF5",X"FFFEF9",X"F5FFFD",X"FFFEFB",X"FCFAFB",X"F8FAF9",X"FFFFFF",X"FFFFFD",X"FFFFFF",X"F9FEFF",X"F8FFFF",X"FFF9ED",X"FFFFF8",X"FCFFFF",X"F7F7F9",X"F8FFFE",X"F0FFFF",X"F7FFFF",X"FFF9FF",X"EBF8FF",X"F8FDFF",X"FFFFFB",X"FFFEFB",X"FCFCFC",X"FCFDFF",X"FCFCFC",X"FFFFFB",X"FEFFFF",X"F9F3F7",X"FFFCFF",X"F8FFFF",X"F6FFFF",X"FFFEFF",X"FFFEFB",X"FBFFF8",X"FFFCF9",X"FFFDFE",X"FFF9FF",X"FFF9FF",X"FFFCF9",X"FEFFFA",X"FCFFFF",X"FBFCFF",X"FFFCFA",X"FFFBFF",X"F7F0F8",X"FFFDFF",X"FFFFFF",X"FDFEFF",X"FAFDFF",X"F8FCFF",X"FFF7FE",X"FBFFFF",X"F2FCFB",X"F9F9F7",X"FFFFFA",X"F7FFFA",X"FBFFFF",X"FFFAFF",X"F2FFFF",X"FFFEFF",X"FFF5FC",X"FFFAFF",X"FAFBFF",X"F8FFFF",X"F6FFFA",X"FFFFF8",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FEFEFE",X"F8FFFF",X"FCFFFF",X"FEFFFD",X"F2FCF3",X"F4FFFA",X"F4FFFF",X"EEF6F8",X"FFFEFF",X"F5FFFF",X"F9FFFF",X"FCFFFF",X"FCFFFF",X"F4FDFC",X"F3FDFC",X"FCFFFF",X"FFFFFB",X"FFFAFC",X"FCFCFE",X"FCFFFF",X"FDFFFC",X"FFFFFA",X"FFFFFB",X"F5F9FC",X"F5FEFF",X"FFFEF6",X"FFFDF4",X"FFFEF3",X"FFFDF6",X"FDFEFF",X"FEFEFF",X"FFF8FF",X"FFF6FF",X"FEFFFF",X"FEFFFF",X"FFFBFF",X"FFF6FF",X"FFF9FF",X"FFFAFF",X"FFFDFF",X"FAFDFF",X"FFFCFD",X"FEFCFD",X"FFFFFF",X"FFFFFF",X"FAFAFC",X"F8F8FA",X"FFFEFF",X"FFFEFF",X"F2FEFE",X"FCFCFF",X"FFF8FF",X"FFFBFF",X"FFFFFF",X"FCFFFB",X"FEFDFB",X"FFF6FD",X"FFFEFA",X"FFF9FD",X"FFFBFF",X"FFFAFF",X"FFFEFF",X"FFFEFF",X"FEF4FC",X"FFF9FF",X"F5FFFF",X"EEF5EE",X"FFFFF8",X"FEF9F6",X"FFFEFF",X"F8F8FF",X"FFFEFF",X"FFFDFF",X"FFFAFA",X"FFF3F3",X"FFFDFD",X"FFFDFE",X"FFFFFF",X"FFFEFF",X"FFFAFC",X"FFFAFB",X"FEFEFF",X"FEFEFF",X"FEFEFF",X"FEFEFF",X"FEFEFF",X"FEFEFF",X"FEFDFF",X"FEFDFF",X"F0FFFD",X"FFFBFF",X"F9FFFF",X"E6FBF2",X"FFFCF6",X"FFF8F8",X"FEF7FE",X"FAF9FF",X"F6FAFD",X"F8FEFE",X"F9FFFF",X"FBFFFF",X"F4F3F8",X"FDFCFF",X"FBFFFF",X"F4FFFE",X"F6FBFF",X"FFFEFF",X"FFFAFF",X"FFF8FF",X"FFF9FC",X"FFFEFD",X"FFFEFF",X"FFF8FF",X"FDF4FF",X"FFFDFF",X"F7FDF9",X"FCFFF6",X"FDFDF5",X"FFFCF9",X"FFFDFB",X"FEF6F3",X"FBFBFD",X"F5F9FA",X"F9FFFF",X"F9FFFF",X"F9FDFC",X"FEFFFF",X"F4F9FC",X"F9FFFF",X"EEFDF6",X"FBFFFA",X"FEFDF8",X"FBFAF8",X"FFFFFF",X"FCFCFA",X"FFFFF4",X"FFFEEB",X"F2FFFD",X"F4FDF8",X"FBFAF6",X"FFFCFC",X"FEFCFD",X"FAFEFF",X"FDFDFF",X"FEFCFF",X"FFFFF8",X"F8F8F0"),
(X"FAF5F2",X"F8F2FE",X"E2EEFF",X"D4FEFF",X"D0FFFF",X"DDF2FF",X"EEF4FF",X"E1EBEA",X"DCEFEB",X"E9FEF9",X"DDF2ED",X"DFEFEC",X"FBFFFF",X"F8F6F9",X"FFFDFF",X"F9F7FA",X"FCD9FF",X"FCCAFF",X"FFD8FF",X"FFD2FF",X"FFE0FF",X"FFDFFF",X"FFDAFF",X"FFCDFF",X"FFCAFF",X"FFC2F8",X"FFE9FF",X"FDF8FF",X"F6FCFC",X"F6FFFF",X"E2FFF8",X"D0FFF6",X"8FFFF1",X"8EFFF0",X"91FFEF",X"A5FFF2",X"C3FFF5",X"D1EEE9",X"E8EDF0",X"E5E3E8",X"FFD6FF",X"FFD1FF",X"FFE5FF",X"FFF2FF",X"FFF5FF",X"FFFDFF",X"FFFDFF",X"FAF3FF",X"FEFFFF",X"FCFFFF",X"F6F7FC",X"FFFDFB",X"FFF1FC",X"F9CCF7",X"FFD2FF",X"FFC9FF",X"EDE4F7",X"F8EFFF",X"E2EDF3",X"BEFBEC",X"ABFFF5",X"A2FFEB",X"C0FEE7",X"F4FFFA",X"F9FFFA",X"F7FFFA",X"F7FFFB",X"E8FFF9",X"B8FFEA",X"9BFFF4",X"87FFED",X"92FFF0",X"8EFFED",X"B6FFF9",X"B5FFF3",X"B5FFF3",X"CCFFFC",X"DDFFFF",X"EBFFFF",X"FDF3FC",X"FDFDFB",X"FFFAFA",X"FFF9FA",X"FFFCFF",X"FFFEFF",X"FEFFFF",X"FBFFFE",X"FDFFFE",X"FFFEFF",X"FBFCFF",X"FFFFF8",X"FFF6E6",X"FADFCE",X"FFF2E6",X"FAF5F1",X"F4FFFF",X"FFFEFF",X"FDFBFC",X"FEFCFD",X"FFFEFF",X"FFFCFF",X"FFFCFF",X"FEF8FC",X"F4EEF2",X"FFD5E8",X"FFCDE6",X"FCE5F7",X"E3EDEC",X"F3F3EB",X"FAEDE4",X"FCF9F2",X"FEFFFF",X"FFFEFB",X"FFFFFD",X"FEFFFF",X"FEFFFF",X"F4F5F7",X"FCFFFF",X"DEE8F2",X"DAEAFA",X"C0F6FF",X"A8F2FF",X"B6FDFF",X"C8F4FF",X"C7EFFF",X"B7F1FF",X"BBF6FF",X"BFE8FF",X"E4F6FF",X"F9FFFF",X"FEFAF7",X"FFFBF7",X"F9F9FB",X"FBFFFF",X"FEFFFF",X"FFFBF8",X"FFF8FF",X"FFFAFF",X"FEFEFF",X"FAFEFF",X"F7F6FB",X"F9E2E8",X"FFD1DB",X"FFC7D5",X"FFC6CC",X"FFC8D1",X"FFC8D9",X"FFCFE5",X"FFC5D5",X"FFC9D5",X"FFC9D9",X"FFCDE5",X"FFDADF",X"FFF0F6",X"FFFCFF",X"F7FFFA",X"EFFFF1",X"F1FFF0",X"FFFFFF",X"FFF8FF",X"FFF9FF",X"FCFFFF",X"FBFFFF",X"FFFEFD",X"E9F0E8",X"D7EDE1",X"E4E2E7",X"FFD5EF",X"FFC3FE",X"FFC9F9",X"FFC5F2",X"FFC9FA",X"FFC2F7",X"FFBBEF",X"FFE6FF",X"FFF3FD",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"F9FAFC",X"FDFBFE",X"F5F3F8",X"DDE1EA",X"DDF7FF",X"C6FAFF",X"B2FFFF",X"A4FFFF",X"BDF5FF",X"E1FFFF",X"F3FDFE",X"FCF6F8",X"FFF8FD",X"FFFDFF",X"FFFEFF",X"FEF9F3",X"FFFEFF",X"FEFEFF",X"FCFFFF",X"F8F8F6",X"FFFEFB",X"FFFFFF",X"EFFCFF",X"E9FFFF",X"BDFAFF",X"D1F8FF",X"EFFDFD",X"FFFDF4",X"FFFCF5",X"FBFFFC",X"F8FFFF",X"F6FFFF",X"FFFEF5",X"F1F1EF",X"F2E9EE",X"FFDDE6",X"FFCBD6",X"FFC9D6",X"FFD4E1",X"FFDAE7",X"FBF7F8",X"FEFCFD",X"FCFAFB",X"FFFFFF",X"FFFFFF",X"FAFAFC",X"F9F9FB",X"EAE8EB",X"FFD9FA",X"FFBFF2",X"FFC1F9",X"FFD2F5",X"EEDFE6",X"FDFEF8",X"FFFEFD",X"FFFAFF",X"FFF8FF",X"FFEDFF",X"FFECFF",X"FFD7F6",X"FFCCEC",X"FFCEEA",X"F0D3E5",X"D0E2E6",X"DAE8FF",X"EEF3FF",X"FFFCFF",X"F9F3F3",X"FFFFFD",X"F9FDFE",X"FFFEFF",X"FFFBFF",X"FFF1F0",X"FFFFFB",X"EEFFFC",X"E4FFFC",X"D5F6EF",X"E5FAF5",X"FEFFFF",X"FFF7FB",X"FEFEFE",X"FEFEFF",X"FEFEFF",X"FEFEFF",X"FDFDFF",X"FDFCFF",X"FCFBFF",X"FCFBFF",X"FFD7FF",X"FFC9FF",X"FFE4FF",X"FFFCFF",X"FFF9FF",X"FFF8F5",X"FCFDF7",X"F7FFFF",X"FFFBFF",X"FFFEFF",X"F2F4F1",X"FEFFFA",X"FEFFFF",X"E7EFFF",X"D0E6FF",X"C6E8FF",X"C1F5FF",X"C7EDFF",X"DCEEFC",X"F7FBFF",X"F4F9FD",X"F8FEFA",X"F3F8F2",X"FFFEFF",X"EAEDFF",X"DBE4F3",X"F1FFFC",X"EAFCEE",X"F7FFFB",X"FCFCFF",X"F9F7FF",X"FFFDFF",X"FFFDFA",X"FFFEFB",X"FAFCF9",X"F7F9F8",X"F3F3F5",X"EDEAF1",X"E2E2EA",X"E6EBF1",X"F0E3F7",X"F0E4F0",X"FBF1F9",X"F8F8FA",X"FEFFFF",X"FFFAF0",X"FFF0D8",X"FFDDB8",X"FFD396",X"FFE1A9",X"FFD39C",X"FFD89D",X"FFE8B5",X"FFE1C4",X"EFDBD4",X"ECECEE",X"E7E7DF",X"FEFEF6"),
(X"F3EEEB",X"B2ACB8",X"6F7B91",X"547E94",X"6998AC",X"768BA0",X"404652",X"000605",X"000602",X"647974",X"455A55",X"485855",X"F0F6F6",X"FBF9FC",X"FDF8FC",X"DAD8DB",X"3C1943",X"45134E",X"43064C",X"3F0748",X"3A1040",X"3A1741",X"43144B",X"4B0E54",X"60155A",X"59184E",X"E5BEDB",X"FEF9FF",X"F4FAFA",X"F8FFFF",X"CFEDE5",X"70A696",X"29B68B",X"2EBB90",X"2BB289",X"43B090",X"3F8471",X"001510",X"000104",X"0A080D",X"430C4F",X"5A2961",X"B188B2",X"D1B7D0",X"DFD4E2",X"FAF8FF",X"FFFDFF",X"FFFBFF",X"F9FAFC",X"F5F8FF",X"FEFFFF",X"FFFDFB",X"E0C6D1",X"481B46",X"5A206A",X"5B1B71",X"20172A",X"04000C",X"000309",X"306D5E",X"49B593",X"42B08B",X"6FAD96",X"E7F4ED",X"F6FFF7",X"F1FEF4",X"F2FFF6",X"C5DFD6",X"559D87",X"29A782",X"2AB890",X"3CBE9A",X"2EB28D",X"48A18B",X"429380",X"63B8A1",X"99D9C9",X"B3E2D8",X"DBF8F4",X"FFFBFF",X"FFFFFD",X"FFFAFA",X"FFF9FA",X"FFFCFF",X"FFFEFF",X"FEFFFF",X"FBFFFE",X"FEFFFF",X"FDFCFF",X"F6F7FB",X"FFFFF8",X"F2E5D5",X"220700",X"FFE7DB",X"FFFEFA",X"F3FFFF",X"FFFEFF",X"FFFDFE",X"FFFEFF",X"FFFCFD",X"FEF9FD",X"FFF9FD",X"F9F3F7",X"EEE8EC",X"8D5C6F",X"430B24",X"0E0009",X"000302",X"65655D",X"D7CAC1",X"F5F2EB",X"FDFFFE",X"FFFEFB",X"FCFBF9",X"FAFBFD",X"FEFFFF",X"FEFFFF",X"F6F9FE",X"96A0AA",X"2C3C4C",X"2C6290",X"206A99",X"175E96",X"224E8B",X"1F477B",X"215B83",X"27628E",X"1A437B",X"95A7B5",X"EEF5FB",X"FFFCF9",X"FFFEFA",X"FCFCFE",X"FAFFFF",X"FCFDFF",X"FFFEFB",X"FFFBFF",X"FFFDFF",X"F0F0F2",X"FCFFFF",X"FFFEFF",X"9B848A",X"591721",X"77111F",X"7F1016",X"751A23",X"611021",X"5D051B",X"6E1020",X"6D131F",X"610919",X"73142C",X"83565B",X"A8898F",X"C3BABD",X"E7F2EA",X"F1FFF3",X"F7FFF6",X"FBFBFB",X"FFF9FF",X"FFFBFF",X"F7FBFC",X"F9FFFF",X"F8F4F3",X"AAB1A9",X"374D41",X"0A080D",X"2B0017",X"740C47",X"661444",X"721B48",X"6A0E3F",X"7C1449",X"781448",X"E5B9D4",X"FFF5FF",X"FDFDFD",X"FDFDFD",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFFFF",X"FEFCFF",X"DBD9DE",X"02060F",X"233D4C",X"578BA3",X"3483A4",X"2F8FB5",X"397180",X"B6D8E1",X"F8FFFF",X"FFFDFF",X"FFFCFF",X"FCF7FD",X"FFFBFC",X"FFFEF8",X"FFFEFF",X"FFFFFF",X"FBFFFE",X"FAFAF8",X"FFFEFB",X"FBFBFB",X"F3FFFF",X"D8F3FC",X"387594",X"CAF1FF",X"F5FFFF",X"FEFBF2",X"FFFFF8",X"FCFFFD",X"F2FCFB",X"F7FFFF",X"FFFEF5",X"FFFFFD",X"A69DA2",X"2F0710",X"5F1621",X"620C19",X"5B1724",X"2E000D",X"D8D4D5",X"FEFCFD",X"FFFEFF",X"F6F6F6",X"FBFBFD",X"FFFFFF",X"F6F6F8",X"B3B1B4",X"3F0223",X"7C1B4E",X"80174F",X"59193C",X"9B8C93",X"F7F8F2",X"FFFDFC",X"F7F2F8",X"FFFBFF",X"FFF0FF",X"E3BBD6",X"93607F",X"571636",X"510F2B",X"120007",X"000509",X"0B1956",X"ABB0DA",X"F5F1FF",X"FFFAFA",X"FFFFFD",X"F6FAFB",X"FFFEFF",X"FFFDFF",X"FFFBFA",X"FFFFFB",X"EFFFFD",X"C7E8DF",X"60817A",X"D5EAE5",X"F7F9F8",X"FFF8FC",X"FEFEFE",X"FEFEFF",X"FEFEFF",X"FEFEFF",X"FEFEFF",X"FDFCFF",X"FCFBFF",X"FBFAFF",X"FAC1F4",X"812566",X"E9BFED",X"FAF7FF",X"FFF5FB",X"FFFBF8",X"F9FAF4",X"F4FFFE",X"FFFBFF",X"FFFBFC",X"FEFFFD",X"FDFFF9",X"FBFDFC",X"98A0B3",X"000F40",X"13357C",X"1D518D",X"11375B",X"788A98",X"EFF3FC",X"FBFFFF",X"FBFFFD",X"FAFFF9",X"FEFCFF",X"878AAD",X"313A49",X"D7E8E2",X"F4FFF8",X"F7FFFB",X"FEFEFF",X"FFFDFF",X"FDFBFF",X"FFF8F5",X"FFFDFA",X"FEFFFD",X"FEFFFF",X"CCCCCE",X"050209",X"090911",X"000107",X"07000E",X"281C28",X"D9CFD7",X"FFFFFF",X"F5F7F6",X"FFFEF4",X"D0B49C",X"916540",X"B27235",X"BD642C",X"C6652E",X"AC6429",X"A2703D",X"7A5538",X"130000",X"000002",X"5B5B53",X"E4E4DC"),
(X"FFFDFF",X"FEFEFE",X"ADDBF5",X"016BA9",X"005F9D",X"8CBDDB",X"D0D5D9",X"C6C5CB",X"93A8A3",X"89A29C",X"6A857E",X"4A615B",X"ECFBF8",X"F8FFFF",X"FBFFFF",X"F5FBFB",X"F2CFF7",X"AD62B7",X"770485",X"82138C",X"803786",X"D3AAD6",X"E1BAE7",X"AE7AB8",X"671C71",X"510E53",X"F2C9F1",X"FFFAFF",X"FFFEFF",X"FFFBFF",X"EDF9F7",X"CBF4E6",X"47D0A6",X"18DEA0",X"06D493",X"5FDDB7",X"CCEDE6",X"CCC5CC",X"B3A2AC",X"A18291",X"A16AAB",X"682C6C",X"460442",X"44083B",X"704561",X"AC9899",X"E7E5CE",X"FCFFDC",X"FFF9F7",X"FFFDFF",X"F9FAFF",X"FEFBF4",X"FFF8FE",X"E0B4E7",X"490A63",X"601981",X"00000B",X"AFA1B0",X"DBCFD9",X"BAD9D3",X"7FD8BC",X"40AC88",X"85D0B9",X"DEFFF6",X"FFFEFB",X"FEFFFD",X"FFFEFF",X"F5FFFE",X"9EF8DE",X"0FCB91",X"13E9A9",X"08BD88",X"7FE6CB",X"D7F1F0",X"BCDBD6",X"62C0A6",X"20AF84",X"04C286",X"5AF3C4",X"DEFFFA",X"F8FFFF",X"FBFFFE",X"FFFDFE",X"FFFDFF",X"FFFEFF",X"FEFEFE",X"FEFEFE",X"FFFEFF",X"FFFEFF",X"FCFFFF",X"F9F3F3",X"CCAA8F",X"BA7B45",X"EDAF76",X"FFF8D8",X"FAFFF9",X"FEFDFB",X"FFFDFE",X"FFFEFF",X"FFFEFF",X"FDFBFE",X"FFFDFF",X"FDFBFE",X"F7F2F8",X"F8C6E1",X"AF487D",X"600A3B",X"0E000B",X"6D6966",X"F4EAE1",X"FFFBF9",X"FFFDFF",X"FFFEFF",X"FFFFFF",X"FEFFFF",X"F7F8FA",X"F7F7F7",X"FEFFFF",X"F5F9FF",X"9CA5B4",X"1653BD",X"277DD0",X"12639B",X"86A8CE",X"C3CFE7",X"8FAFC8",X"5386B5",X"1C4795",X"96ABBE",X"F8FFFF",X"FEFAF7",X"FCF7F4",X"FEFFFF",X"FBFFFF",X"FCFDFF",X"FFFDFA",X"FBF6FD",X"FEFFFF",X"FFFFFD",X"FFF7FE",X"FFF8FF",X"FEE4ED",X"F091A5",X"A6001D",X"B4000B",X"BC4A52",X"FCCDD3",X"EED8DB",X"BD9F9F",X"B78787",X"C07884",X"93304C",X"31040B",X"1A0002",X"020100",X"7D947A",X"D1F0C6",X"E9FFDA",X"FBFFF0",X"FFFCFD",X"FFFEFF",X"FBFFFF",X"FDFDFF",X"FFF7F8",X"E4EEE6",X"586D66",X"12000A",X"701040",X"A6276A",X"C182AD",X"D1A8C8",X"B78EAE",X"BB6896",X"791748",X"D8BFD2",X"F0FFFF",X"FDFDFD",X"FDFDFD",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FCF6F6",X"FFFEFD",X"FFFEFF",X"D8DAE6",X"4D5D76",X"25557B",X"449FCC",X"1690C1",X"8AC3CE",X"DEFFFF",X"FAFFFB",X"FFF5F3",X"FFFBFF",X"FFFDFF",X"FFFEFF",X"FFFCF9",X"FDFBFC",X"FEFFFF",X"FCFEFD",X"FFFEFD",X"FFFCFD",X"F7F6FB",X"EEFFFF",X"A6D2DD",X"0484B3",X"6BC4E4",X"D7FBFF",X"FDFBFE",X"FFF8FB",X"FFF8FC",X"FFFEFD",X"FFFFFB",X"FFFCF3",X"FAFBF3",X"F5EDEA",X"A97174",X"7D0B13",X"A01927",X"690310",X"DEA0AB",X"FFFEFD",X"FFFEFF",X"F7F5F6",X"FEFEFE",X"FCFDFF",X"F7F7F9",X"FFFFFF",X"F5F4F9",X"E473AB",X"B5055A",X"B7005B",X"C55C94",X"F1DBE7",X"FFFFFA",X"FCFBF9",X"FAFFFF",X"F9F1FF",X"FF9ACE",X"9B0042",X"952057",X"BB8FA8",X"D3C7D1",X"B7B8BD",X"556769",X"162D79",X"B6C0F5",X"FFFCFF",X"FFFCFB",X"FDFFF9",X"F9FFF9",X"FFFFFA",X"FEF9F3",X"FCFFFD",X"F1FBFA",X"F1FFFF",X"94A9AC",X"051A1D",X"9EABB1",X"FCFFFF",X"FDFAFF",X"FFFFFD",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFF",X"FDFCFF",X"FCFBFF",X"FBFAFF",X"F5B3F3",X"AF0172",X"CE2DA1",X"FFB1FF",X"FFDEFF",X"FCFBFF",X"FEFFFD",X"FFFCFD",X"FFF7F7",X"FFF7FD",X"FFF8FF",X"FFF8F6",X"FFFCFB",X"FAFAFF",X"8A9CE6",X"0D2E9F",X"0044B3",X"77A9E6",X"E5FCFF",X"F4F8FF",X"F7FAFF",X"F5FDFF",X"F2F7FA",X"FEFEFF",X"8D92CC",X"05092F",X"545365",X"F3E9F4",X"FFF7FF",X"FFF0FF",X"FFFBFF",X"FFFFF8",X"FFFEFB",X"FFFEFC",X"F7F7F7",X"FFFEFF",X"F5EFF3",X"E2DCE0",X"6E6C71",X"020307",X"080413",X"B2ADB4",X"FFFAFE",X"FCFDFF",X"FBFFFF",X"FFFAF7",X"FFF2DE",X"E5B08E",X"D25803",X"FA621F",X"E55D21",X"E39D61",X"DFC18F",X"DBBDA5",X"93807A",X"000400",X"31322D",X"E5E6E1"),
(X"FDF7F9",X"FAFAFA",X"BBE9FF",X"0E78B6",X"0771AF",X"B1E2FF",X"FAFFFF",X"FFFEFF",X"F1FFFF",X"E5FEF8",X"CBE6DF",X"79908A",X"F0FFFC",X"F8FFFF",X"F1F7F7",X"F6FCFC",X"FFF0FF",X"CB80D5",X"790687",X"70017A",X"D58CDB",X"FFE2FF",X"FFE3FF",X"FFE4FF",X"FFB6FF",X"9C599E",X"FAD1F9",X"FFFAFF",X"FAF8FD",X"FBF6FA",X"F7FFFF",X"E0FFFB",X"79FFD8",X"0CD294",X"00CA89",X"79F7D1",X"E9FFFF",X"FFF9FF",X"FFF7FF",X"FFEBFA",X"FFDEFF",X"FABEFE",X"E09EDC",X"64285B",X"1F0010",X"100000",X"4A4831",X"E3E9C3",X"FFFDFB",X"FFFCFF",X"FEFFFF",X"F5F2EB",X"FFF9FF",X"FFE7FF",X"A667C0",X"400061",X"555964",X"EBDDEC",X"FFFAFF",X"E2FFFB",X"C4FFFF",X"92FEDA",X"7EC9B2",X"E8FFFF",X"FEF9F6",X"FDFFFC",X"FBF9FA",X"F4FEFD",X"B1FFF1",X"0FCB91",X"02D898",X"2CE1AC",X"A7FFF3",X"EAFFFF",X"E3FFFD",X"B2FFF6",X"67F6CB",X"03C185",X"22BB8C",X"ADD0C9",X"F4FFFB",X"FBFFFE",X"FFFEFF",X"FFFCFE",X"FEFCFD",X"FEFEFE",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"F4F7FE",X"F9F3F3",X"937156",X"CC8D57",X"E4A66D",X"FFE9C9",X"FCFFFB",X"FEFDFB",X"FEFCFD",X"FFFEFF",X"FFFEFF",X"FDFBFE",X"FFFDFF",X"FFFEFF",X"FFFBFF",X"FFE2FD",X"CD669B",X"6A1445",X"0E000B",X"797572",X"FFFAF1",X"FFFCFA",X"FFFCFF",X"FFFCFD",X"FDFDFF",X"FEFFFF",X"FEFFFF",X"FCFCFC",X"F7F8FC",X"FBFFFF",X"B1BAC9",X"002A94",X"247ACD",X"499AD2",X"D5F7FF",X"F2FEFF",X"E0FFFF",X"D2FFFF",X"5580CE",X"879CAF",X"F1FAFF",X"FFFEFB",X"FFFCF9",X"FEFFFF",X"F9FEFF",X"F9FAFE",X"FFFEFB",X"FFFCFF",X"FEFFFF",X"FFFFFD",X"FBEEF5",X"FFF7FF",X"FFF6FF",X"FFB6CA",X"B4092B",X"B8020F",X"D4626A",X"FFE7ED",X"FFF5F8",X"FFEFEF",X"FFE6E6",X"FFDFEB",X"FFB3CF",X"DAADB4",X"694C51",X"010000",X"7F967C",X"708F65",X"B2CBA3",X"FCFFF1",X"FBF2F3",X"FDFBFC",X"FBFFFF",X"FFFFFF",X"FFFCFD",X"F8FFFA",X"71867F",X"0F0007",X"650535",X"CB4C8F",X"FFD5FF",X"FFECFF",X"FFE5FF",X"FFCAF8",X"CF6D9E",X"DEC5D8",X"EFFFFF",X"FDFDFD",X"FDFDFD",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFDFD",X"F7F3F2",X"F8F6F9",X"F9FBFF",X"76869F",X"000C32",X"1F7AA7",X"2BA5D6",X"C5FEFF",X"E4FFFF",X"F9FEFA",X"FFFCFA",X"FFFAFE",X"FDFAFF",X"FFFEFF",X"FFFDFA",X"FEFCFD",X"FEFFFF",X"FAFCFB",X"FFFEFD",X"FFFBFC",X"FFFEFF",X"E7FEFF",X"7AA6B1",X"0989B8",X"48A1C1",X"DCFFFF",X"FEFCFF",X"FFFAFD",X"FFFBFF",X"FCF8F7",X"FDFEF9",X"FFFAF1",X"FFFFF8",X"FFF8F5",X"FFDADD",X"6C0002",X"930C1A",X"87212E",X"FFDDE8",X"F9F5F4",X"FFFEFF",X"FEFCFD",X"FEFEFE",X"F8F9FB",X"FAFAFC",X"FFFFFF",X"F9F8FD",X"FF9CD4",X"B30358",X"B7005B",X"F087BF",X"FFF7FF",X"FCFDF7",X"F6F5F3",X"FBFFFF",X"F6EEFD",X"92275B",X"AB0652",X"FF8AC1",X"FFE8FF",X"FFF8FF",X"F0F1F6",X"E8FAFC",X"536AB6",X"A0AADF",X"FDFAFF",X"FCF8F7",X"F9FCF5",X"F3FAF3",X"FEFFF9",X"FFFEF8",X"F5FAF6",X"F5FFFE",X"E4F6F6",X"263B3E",X"000D10",X"233036",X"E4E7EE",X"FFFDFF",X"FEFEFC",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFF",X"FDFCFF",X"FCFBFF",X"FBFAFF",X"F7B5F5",X"BD0F80",X"EF4EC2",X"AF4BA1",X"F6C0F1",X"FBFAFF",X"F1F3F0",X"FFFBFC",X"FFFAFA",X"FFFBFF",X"FFFCFF",X"FFFDFB",X"FFFBFA",X"FCFCFF",X"B9CBFF",X"3F60D1",X"084CBB",X"75A7E4",X"EAFFFF",X"FBFFFF",X"F6F9FF",X"F4FCFF",X"FBFFFF",X"F8F8FF",X"8F94CE",X"00042A",X"000010",X"776D78",X"F7E5F5",X"FFF8FF",X"FCF1F7",X"FFFFF7",X"FEFAF7",X"FFFFFD",X"FFFFFF",X"FCFAFB",X"FFFAFE",X"FFFDFF",X"AAA8AD",X"000004",X"01000C",X"C0BBC2",X"FFFDFF",X"FAFBFF",X"F4F9FD",X"FFFCF9",X"FFF8E4",X"FDC8A6",X"D35904",X"F65E1B",X"D1490D",X"FFD498",X"FFFCCA",X"FFEAD2",X"FFF4EE",X"8E9A96",X"979893",X"FFFFFB"),
(X"FDFEFF",X"FFFFF6",X"C3E9FF",X"0A6EE0",X"0063D8",X"B6D7FF",X"FFF7F8",X"FCF6FF",X"FFFAFE",X"FEFEFF",X"F8FCFD",X"D9DDDE",X"FFFEFF",X"FCF6FA",X"FFFCFF",X"FFFDFF",X"FBFFF6",X"D29BD4",X"7A0681",X"7C0980",X"DA9FD7",X"FFFCF7",X"F7FFF2",X"F8FDF7",X"FFF0FF",X"DFDFE7",X"F5FFFA",X"F7FDEF",X"FFFEF5",X"FFFFFD",X"F9FFFF",X"F1F9FC",X"B5E7DB",X"1DCA94",X"01DA95",X"87F4D4",X"F9FAFE",X"FEF4FC",X"F7FFFF",X"FAFFFF",X"FFFFF4",X"FFF8FF",X"FFF4FF",X"E4CDEA",X"675257",X"291600",X"A59035",X"D7BF43",X"FEF5B4",X"FCF7DA",X"FCFFFF",X"F9FFFF",X"FEFFFF",X"F8EAFF",X"907890",X"110000",X"796F77",X"F8F9FD",X"F5FFFF",X"F7FFFF",X"EDEFEE",X"F9F7FC",X"E8EBF0",X"F3FEFF",X"FFFEFF",X"F9FDFF",X"FFF6FF",X"FFF3FF",X"CBFFF9",X"40EBB7",X"05C288",X"57DFB7",X"C3FFF2",X"FDF8FF",X"FCFDFF",X"F0FFFF",X"D5F4EC",X"4ECDA4",X"05C687",X"50D8AA",X"E3FAF4",X"F1FFFD",X"FCFFFF",X"FEFCFF",X"FCFAFB",X"FFFDFE",X"FFFEFF",X"FFFBFD",X"FFFDF6",X"FCFFFF",X"C5BAC2",X"370500",X"F09640",X"E48727",X"FFCB92",X"FFFCF2",X"FFFFFD",X"FCFCFA",X"FEFEFE",X"FFFFFF",X"FCFCFE",X"FBFBFD",X"FEFDFF",X"FCFDFF",X"F7F8FF",X"E984C0",X"B5075E",X"710034",X"A58B94",X"FFFBF5",X"FFFBFC",X"E9FFFF",X"FFFEFF",X"FBFEFF",X"FBFEFF",X"FEFFFF",X"FFFEFD",X"FDF9F8",X"FEFDFF",X"CCCFD6",X"040026",X"274C67",X"7DADC1",X"EEF7FF",X"FFFBFF",X"EBF5ED",X"E7FFFF",X"D6F0FF",X"CFE5FA",X"F8FFFF",X"FFF9F9",X"FDF8F5",X"FEFFFF",X"F9FFFF",X"FEFFFF",X"FFFEFB",X"FFFEFF",X"F3FAF3",X"FDFAF5",X"FFF9FF",X"F9FFFF",X"E8FFFD",X"FFDDDE",X"BD4457",X"A8000B",X"BF5E69",X"FFE3EF",X"FFFBFF",X"FFFBFF",X"FBF9FA",X"FBFFFF",X"FBFBFF",X"FFFFFB",X"DFE6DF",X"A0B7A5",X"769D71",X"6D9E5D",X"608E4D",X"AFD6A7",X"EAFFF0",X"FCFFFF",X"F3FCFB",X"FFFBFF",X"FFFAFD",X"EFF5F1",X"91A19E",X"2E001C",X"8E094A",X"D075A0",X"FFECFF",X"FBEEF8",X"EFF9FA",X"FFFCFF",X"FED9EA",X"F6EDEE",X"FFFEF8",X"FDFDFD",X"FDFDFD",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FAF5FC",X"FEFFFF",X"FCFFF8",X"FFFBF1",X"BCAAA6",X"080002",X"000915",X"608691",X"E6F9FF",X"F1F9FC",X"FFFEF5",X"FFFFF4",X"F9FFFB",X"F1FFFF",X"F8FFFF",X"FEFFFD",X"FFFFFF",X"FEFFFF",X"FCFEFD",X"FFFDFD",X"FFF9FB",X"FEFFFF",X"B6D2DD",X"2A606C",X"4A6E88",X"293C4A",X"A3A3A5",X"FFFBF8",X"FFFEFF",X"FAFEFF",X"FEFFFF",X"FFFDFA",X"FBF9FE",X"F1FFFF",X"F4FFFF",X"FCD7DF",X"932A3B",X"7E0015",X"8F4053",X"FFE8F7",X"FFFDFD",X"FFFBFA",X"FBF9FA",X"FFFFFF",X"FEFFFF",X"FAFBFD",X"FEFDFF",X"FFFEFF",X"F8AEDF",X"A6065C",X"BC0768",X"FDA4DA",X"F4F3F9",X"F2FCF3",X"FFFEFD",X"FCFDFF",X"FFD3F3",X"79154B",X"B44D84",X"FFDEFE",X"FFF7FF",X"FFF2FF",X"FFF4FF",X"F4FFFF",X"BEE6EE",X"C1D7D5",X"FCFFF6",X"FEFBF2",X"FEFFFF",X"FBFFFF",X"FAF9FF",X"FFF8FB",X"FEFFFF",X"FFF8FF",X"D8BCD2",X"1A000F",X"491D3E",X"16000F",X"AF99AE",X"FFF9FF",X"FDFDFB",X"FEFEFC",X"FEFEFE",X"FFFFFF",X"FEFEFF",X"FDFDFF",X"FBFBFD",X"FBFBFD",X"F0B4E7",X"A50066",X"FF63E9",X"CC32B4",X"DF4DB8",X"FFC5FF",X"FFE6FF",X"FEF7FF",X"F8FFF8",X"F9FFFF",X"EFF2FF",X"FFFEFD",X"FFFEEB",X"F9FBED",X"EAFFFF",X"557CB5",X"0E3DB1",X"9AB5EA",X"FEFFFD",X"FFFCF3",X"FFF8F8",X"FFFEFC",X"FEFFFF",X"F8F9FE",X"87A2B7",X"000310",X"3D3A45",X"180014",X"946F91",X"FFE6FF",X"FFFAFF",X"F3F9F5",X"F8FFFF",X"F4FDFC",X"F5FBFB",X"FEFFFF",X"FEF9FD",X"FFFEFF",X"C5C5C3",X"0C130C",X"1A3B2A",X"CDE2D1",X"F8FEF4",X"FEFFFF",X"FBFFFF",X"FBF9FF",X"FFF5F1",X"F5D6C2",X"DC6D13",X"E65B20",X"E67E5B",X"F4E3C7",X"EEFFF2",X"FFF9FE",X"FFEEF4",X"FFFAF5",X"E0E0E2",X"FBFBFD"),
(X"F9FAFC",X"FFFFF6",X"C0E6FF",X"1377E9",X"096CE1",X"B4D5FF",X"FFFBFC",X"FFFCFF",X"FFFAFE",X"FEFEFF",X"FBFFFF",X"FCFFFF",X"FDFBFE",X"FFFDFF",X"FFFCFF",X"FEF8FC",X"F4FCEF",X"F3BCF5",X"700077",X"6D0071",X"ECB1E9",X"FEFBF6",X"F8FFF3",X"F9FEF8",X"FFF2FF",X"FEFEFF",X"EEFEF3",X"FCFFF4",X"FFFFF6",X"F6F6F4",X"F6FEFF",X"F9FFFF",X"BDEFE3",X"27D49E",X"00D994",X"7EEBCB",X"FEFFFF",X"FFFBFF",X"F2FEFE",X"FAFFFF",X"FBFBEF",X"FFFBFF",X"FFF4FF",X"FFF2FF",X"EFDADF",X"B7A47A",X"CFBA5F",X"C8B034",X"E2D998",X"FFFDE0",X"F8FCFB",X"F1F9FB",X"FAFBFF",X"FFF7FF",X"9D859D",X"120001",X"7A7078",X"FAFBFF",X"F3FFFD",X"F5FFFD",X"FEFFFF",X"FCFAFF",X"F7FAFF",X"F7FFFF",X"FDFBFF",X"FBFFFF",X"FFF9FF",X"FFF0FD",X"CAFFF8",X"40EBB7",X"15D298",X"4CD4AC",X"C8FFF7",X"FFFBFF",X"FBFCFF",X"EEFFFF",X"E3FFFA",X"6DECC3",X"0DCE8F",X"3FC799",X"DBF2EC",X"EEFDFA",X"FCFFFF",X"FDFBFE",X"FBF9FA",X"FFFDFE",X"FFFEFF",X"FFF9FB",X"FCF9F2",X"FCFFFF",X"8E838B",X"5F2D0C",X"F09640",X"E18424",X"DEAA71",X"FEF4EA",X"FFFFFD",X"FAFAF8",X"FCFCFC",X"FFFFFF",X"FEFEFF",X"FCFCFE",X"FFFEFF",X"FEFFFF",X"F7F8FF",X"F994D0",X"B90B62",X"8B144E",X"BAA0A9",X"FFF8F2",X"FFFCFD",X"EEFFFF",X"FEFDFF",X"FCFFFF",X"FCFFFF",X"FBFCFE",X"FFFDFC",X"FFFEFD",X"FAF9FE",X"E2E5EC",X"48416A",X"000823",X"76A6BA",X"F0F9FF",X"FFF9FD",X"F9FFFB",X"E1FFFF",X"EBFFFF",X"EAFFFF",X"F7FFFF",X"FDF7F7",X"FFFEFB",X"FEFFFF",X"F6FDFF",X"FEFFFF",X"FFFBF8",X"FFFDFE",X"FBFFFB",X"FFFEF9",X"FFF5FB",X"F7FFFF",X"ECFFFF",X"FFE6E7",X"CA5164",X"A7000A",X"C2616C",X"FADEEA",X"FFFBFF",X"FFF9FF",X"FFFEFF",X"FAFEFF",X"FEFEFF",X"FAF9F5",X"FBFFFB",X"EBFFF0",X"A4CB9F",X"659655",X"709E5D",X"688F60",X"C2E3C8",X"FAFEFD",X"F7FFFF",X"FCF7FB",X"FFFAFD",X"F9FFFB",X"A6B6B3",X"21000F",X"840040",X"DC81AC",X"FFE8FC",X"FFFAFF",X"F7FFFF",X"FDF6FE",X"FFF2FF",X"FFFCFD",X"FFFBF5",X"FDFDFD",X"FEFEFE",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFDFF",X"FAFCFB",X"F4FAF0",X"FFFEF4",X"C6B4B0",X"0D0007",X"00020E",X"3F6570",X"E1F4FF",X"F9FFFF",X"FFFFF6",X"FDF9EE",X"FBFFFD",X"F5FFFF",X"F6FFFF",X"FEFFFD",X"FBFBFB",X"FEFFFF",X"FEFFFF",X"FFF9F9",X"FFF7F9",X"FCFDFF",X"77939E",X"000F1B",X"000822",X"000412",X"555557",X"F4EFEC",X"FCFBFF",X"F7FBFF",X"FAFBFF",X"FFFDFA",X"FFFEFF",X"ECFEFF",X"F4FFFF",X"FFE4EC",X"AB4253",X"820419",X"A7586B",X"FFE6F5",X"FFFDFD",X"FCF8F7",X"FEFCFD",X"FEFEFE",X"FCFDFF",X"FDFEFF",X"FDFCFF",X"FEFDFF",X"FFBDEE",X"B9196F",X"B70263",X"FFB0E6",X"FFFEFF",X"F8FFF9",X"FAF6F5",X"FEFFFF",X"FFD3F3",X"69053B",X"6B043B",X"E2B9D9",X"FFF7FF",X"FFF5FF",X"FFEAF7",X"F1FFFF",X"E0FFFF",X"EDFFFF",X"FEFFF8",X"FFFEF5",X"FCFDFF",X"FAFEFF",X"F8F7FF",X"FFFCFF",X"F5F6FA",X"FFFAFF",X"91758B",X"724967",X"9C7091",X"583651",X"AD97AC",X"F9ECFD",X"FCFCFA",X"FDFDFB",X"FEFEFE",X"FEFEFF",X"FEFEFF",X"FCFCFE",X"FBFBFD",X"FAFAFC",X"F1B5E8",X"B50776",X"B90B91",X"C52BAD",X"A10F7A",X"B25A97",X"FFD5F1",X"FCF5FD",X"F9FFF9",X"F7FEFF",X"FAFDFF",X"FDF9F8",X"FFFCE9",X"FFFFF3",X"E7FDFF",X"5F86BF",X"0130A4",X"ACC7FC",X"FEFFFD",X"FFF8EF",X"FFF8F8",X"FFFFFD",X"FAFCFB",X"FEFFFF",X"849FB4",X"000B18",X"010009",X"240B20",X"3A1537",X"C3A4C4",X"FBF0FE",X"F8FEFA",X"F6FFFE",X"F9FFFF",X"F9FFFF",X"FEFFFF",X"FFFAFE",X"FFFDFE",X"DFDFDD",X"000700",X"355645",X"D2E7D6",X"FBFFF7",X"FEFFFF",X"F4F8FF",X"FFFDFF",X"FFF7F3",X"FBDCC8",X"D6670D",X"DA4F14",X"EB8360",X"FFF6DA",X"F0FFF4",X"FFF6FB",X"FFF1F7",X"FFFDF8",X"FFFFFF",X"FFFFFF"),
(X"FFF3FF",X"FFFDFD",X"BEEEFC",X"0F7BC6",X"0971E0",X"B1E6F6",X"FEFEFF",X"FFFAF7",X"FCFBFF",X"F9FDFF",X"EEF9F5",X"F8FFFC",X"FBFDF8",X"FEFAF9",X"FFF9FB",X"FFFDFF",X"FFFDF7",X"E3C5DD",X"2A0F30",X"140012",X"CAB6BF",X"F7FFFF",X"EEFFF8",X"FFFCF0",X"EEFFFF",X"F5FAFD",X"FFFFFF",X"FFFEFF",X"FFF9FC",X"FEFAFB",X"FDFDFF",X"FFFDFF",X"CFE6DE",X"22D498",X"0FD192",X"8ABDAE",X"FEFEFF",X"FFFDFF",X"FFF4FF",X"ECFFFF",X"FEF9F6",X"FFFDFA",X"FFFDFD",X"FAF8F9",X"FEFCED",X"F3EAA9",X"C3AC2A",X"D6B202",X"C8BD09",X"F5EEA6",X"FFFFEC",X"F5FAFE",X"FEFBFF",X"FFEDFF",X"BC94B6",X"000107",X"7E747D",X"FFF5F9",X"FFF6FD",X"FEFEFF",X"F4FFFF",X"F7FFF7",X"F3FDF4",X"FFFAFF",X"EEFFFD",X"FFF3FC",X"FEFFFF",X"FAFFFF",X"E0FDF8",X"81DEC1",X"31C190",X"69AD94",X"F1FFF2",X"F8FFFA",X"FAFCF9",X"FFFCFF",X"F3FCFF",X"8AB1AE",X"327261",X"72BD9F",X"DEF6FF",X"F5FCFF",X"FFF7FC",X"FFFCF8",X"F0FFF6",X"F5FFFA",X"FFFEFF",X"F1FAF7",X"FFF8FF",X"D2EBF2",X"000209",X"9E7F7A",X"F6C791",X"E08211",X"EE881C",X"FFE4AD",X"F5FDF0",X"FFFDFA",X"FEF9FD",X"FFF9FF",X"FFFAFF",X"FEFFFD",X"EAF9F2",X"FFFEFF",X"FDFDFB",X"EEB4C2",X"D1005C",X"CF0170",X"EBB9D6",X"FFFDFA",X"FFF8FF",X"FCFEF9",X"FFFAFF",X"FFFBFF",X"FDFDFF",X"FEFEFE",X"FFFDFF",X"FFFAFF",X"FDF8FE",X"F5F7E9",X"665B59",X"050100",X"8C8A8D",X"FFFFFD",X"F4F4FC",X"F8FEFF",X"F5FFF3",X"F6FDF6",X"FCFBFF",X"F8F8FA",X"FEFEFC",X"FFFFFB",X"FEFFFA",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FEFEFE",X"FBFFFC",X"F9FFFD",X"FFFDFF",X"FFFAFF",X"F4FFFF",X"FEEEF1",X"C2667D",X"990000",X"A8565C",X"F8DEEB",X"FFF9FF",X"FFF6FA",X"FEFFFF",X"F0FFFF",X"FFFCFD",X"FFFFF7",X"FAF7FE",X"FDFBFF",X"F4FFFB",X"8BA683",X"69945C",X"6C9B67",X"8BB992",X"FAFCEF",X"FFFFFD",X"FCFAFF",X"FFF9FD",X"FEFEF6",X"D3C9C7",X"3A0013",X"99004C",X"E195C4",X"FEFBFF",X"FCFCFF",X"FFFBFF",X"FEFFFF",X"FFFFFF",X"FEFFFF",X"FFF2FF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"F2FFFA",X"FFF0FF",X"FFFAFF",X"F5FDF0",X"DBD3E2",X"0B000E",X"010002",X"687073",X"F2F5FC",X"FFF7FF",X"FFF8FF",X"FDFCFF",X"F8FFFF",X"FCFFFF",X"FDFFFC",X"FBFFF8",X"F8F8FA",X"FBFFFF",X"FFFCFF",X"FEEAF5",X"FFF9FF",X"E9E3E3",X"030002",X"5E4E59",X"9D8D98",X"110001",X"1C0000",X"E5BAC1",X"FFFAFB",X"EEFDFA",X"F3FEFF",X"FFF8FF",X"F9FFF5",X"FFFEFF",X"FBFAFF",X"F9EEF2",X"A2696F",X"640211",X"BA6D7F",X"FFEBF6",X"FFFDFF",X"FDFEFF",X"F8FFFC",X"F8FFFF",X"F9FFFF",X"FCFDFF",X"FEFCFF",X"FFFEFC",X"FFD6F3",X"703C53",X"643C45",X"E8DCDC",X"FDFBFE",X"FFF9FF",X"FFFBFF",X"F4FFF8",X"F0E5ED",X"0E0824",X"00002B",X"34436E",X"DBEDFF",X"F5FFFF",X"F1F5F4",X"FFFEFF",X"FAF9FF",X"F8FFFF",X"F8FFFF",X"FEFEF4",X"FFFFFA",X"F8FFFF",X"F4F6FF",X"FFF9FF",X"FFFDF1",X"DAEFF0",X"3A354C",X"B788B4",X"F4ADF1",X"CE4EBB",X"D649B9",X"FFC1FF",X"FFF5FF",X"F9FFFF",X"F2FFFF",X"F2F6F9",X"FFFDFF",X"FBFFFE",X"F7F7F5",X"FFF7FA",X"FFB4ED",X"A70980",X"F27BDF",X"D277BC",X"B41482",X"C80E95",X"CC48AD",X"FFC9FF",X"FFF3FF",X"FCF9FF",X"FBFAFF",X"FCFCFA",X"F9FFF8",X"FFFCFB",X"FCFBFF",X"6790A6",X"104480",X"B9D1ED",X"FAFFFC",X"FFFFFA",X"FFFFFF",X"F9FBFA",X"FFFEFF",X"FEFFFF",X"8B8796",X"5C4C69",X"928F98",X"03010E",X"CE2CA3",X"E63ECF",X"FF8BF4",X"FFE3FF",X"F3F7FA",X"FFFCFD",X"FFF7F4",X"F5FAF4",X"F9FFFF",X"FAFBFF",X"E7EAF1",X"000606",X"4B5E62",X"E6F5F2",X"FFFBF8",X"FFFAFD",X"FFFBFF",X"F9FFFF",X"FFF6F9",X"FFDEE2",X"CB774B",X"E3490D",X"EE8F63",X"FCFEE9",X"F9F4E1",X"FFFBFC",X"F0FCFF",X"FFF4FB",X"FFFBF5",X"F4F8F7"),
(X"FFF5FF",X"FFFDFD",X"CDFDFF",X"1682CD",X"0870DF",X"A4D9E9",X"FEFEFF",X"FFFAF7",X"FAF9FF",X"FCFFFF",X"F3FEFA",X"F8FFFC",X"FEFFFB",X"F8F4F3",X"FFFDFF",X"F7F1F5",X"FEF9F3",X"ECCEE6",X"17001D",X"0D000B",X"D5C1CA",X"F4FEFD",X"EDFFF7",X"FFF7EB",X"F2FFFF",X"F9FEFF",X"FFFFFF",X"FAF6F7",X"FFFBFE",X"FFFEFF",X"FEFEFF",X"FEFCFF",X"CEE5DD",X"26D89C",X"00B879",X"82B5A6",X"FFFFFF",X"FFFAFE",X"FFF5FF",X"ECFFFF",X"FFFEFB",X"FFFDFA",X"FDF7F7",X"FAF8F9",X"FFFFF1",X"FFFBBA",X"DCC543",X"DAB606",X"C7BC08",X"E1DA92",X"FFFFEA",X"F7FCFF",X"FDFAFF",X"FFF2FF",X"C8A0C2",X"000208",X"756B74",X"FFF4F8",X"FFF8FF",X"F8F8FF",X"F1FFFF",X"F2FEF2",X"F4FEF5",X"FFFDFF",X"EDFFFC",X"FFF6FF",X"FEFFFF",X"F7FCFF",X"E4FFFC",X"89E6C9",X"008150",X"377B62",X"EAF8EB",X"F0FCF2",X"FEFFFD",X"FBF6FC",X"F3FCFF",X"79A09D",X"001706",X"59A486",X"E5FDFF",X"F5FCFF",X"FFF4F9",X"FFF7F3",X"F0FFF6",X"F6FFFB",X"FFFDFE",X"F5FEFB",X"FFF7FE",X"B0C9D0",X"00060D",X"E2C3BE",X"FFD9A3",X"F59726",X"DE780C",X"DEB982",X"FBFFF6",X"FFFCF9",X"FFFDFF",X"FFF8FF",X"FFF5FC",X"FEFFFD",X"F3FFFB",X"FFFEFF",X"FFFFFD",X"EFB5C3",X"D3005E",X"D20473",X"F4C2DF",X"FFFEFB",X"FFF8FF",X"FEFFFB",X"FFFAFF",X"FFFCFF",X"FEFEFF",X"FEFEFE",X"FFFDFF",X"FFFBFF",X"FFFAFF",X"F8FAEC",X"776C6A",X"080400",X"838184",X"FCFBF9",X"FEFEFF",X"F9FFFF",X"F4FFF2",X"FBFFFB",X"FDFCFF",X"FFFFFF",X"FEFEFC",X"FCFDF8",X"FBFCF7",X"FCFCFC",X"FFFEFF",X"FFFEFF",X"FEFEFE",X"FBFFFC",X"FAFFFE",X"FFFDFF",X"FFFBFF",X"F6FFFF",X"FFF2F5",X"C96D84",X"9A0100",X"A45258",X"F7DDEA",X"FFF9FF",X"FFF5F9",X"FEFFFF",X"EFFFFF",X"FFFCFD",X"FFFFF7",X"FFFDFF",X"FCFAFF",X"F5FFFC",X"C2DDBA",X"6A955D",X"6F9E6A",X"6F9D76",X"E2E4D7",X"FFFFFD",X"FFFEFF",X"FEF8FC",X"FFFFF8",X"DCD2D0",X"45001E",X"9C014F",X"ECA0CF",X"F2EFFF",X"FEFEFF",X"FFFCFF",X"FBFDFC",X"FDFDFF",X"FAFBFF",X"FFF7FF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"F0FFF8",X"FFF2FF",X"FFF8FD",X"F9FFF4",X"E5DDEC",X"0B000E",X"010002",X"7F878A",X"F4F7FE",X"FFF8FF",X"FFF8FF",X"FDFCFF",X"F8FFFF",X"FCFFFF",X"FDFFFC",X"FBFFF8",X"FFFFFF",X"F2F7FA",X"FFFDFF",X"FFF0FB",X"FFF9FF",X"A59F9F",X"030002",X"CABAC5",X"E0D0DB",X"1A050A",X"2A060A",X"9F747B",X"FFF1F2",X"F5FFFF",X"F2FDFF",X"FFF5FF",X"F9FFF5",X"FFFDFE",X"FFFEFF",X"FDF2F6",X"B0777D",X"650312",X"C5788A",X"FFF3FE",X"FFFDFF",X"FCFDFF",X"F7FFFB",X"F8FFFF",X"F9FFFF",X"FCFDFF",X"FEFCFF",X"FFFFFD",X"FFD8F5",X"5B273E",X"4A222B",X"E6DADA",X"FFFEFF",X"FFF6FF",X"FDF8FC",X"F7FFFB",X"F7ECF4",X"48425E",X"191D4C",X"071641",X"63758D",X"DAE8EB",X"FCFFFF",X"FBF9FA",X"FFFEFF",X"F6FFFF",X"F4FEFF",X"FFFFF6",X"FEFFF9",X"F0F9FF",X"FCFEFF",X"FFF4FC",X"FFFFF3",X"9EB3B4",X"010013",X"F3C4F0",X"FFCBFF",X"CA4AB7",X"A21585",X"E198DF",X"FFF5FF",X"F4FCFF",X"EAFCFC",X"FCFFFF",X"FFFBFF",X"F9FDFC",X"FFFFFD",X"FFF6F9",X"FFB8F1",X"A00279",X"FF93F7",X"FFCAFF",X"F555C3",X"E127AE",X"C844A9",X"BC67A8",X"F8DAE6",X"F9F6FD",X"FFFEFF",X"FFFFFD",X"F7FFF6",X"FBF7F6",X"FAF9FF",X"5D869C",X"174B87",X"CBE3FF",X"FBFFFD",X"FFFFFA",X"FFFFFF",X"FBFDFC",X"FFFCFD",X"F9FAFF",X"74707F",X"1A0A27",X"F2EFF8",X"AFADBA",X"AE0C83",X"D32BBC",X"9B0C75",X"E3BDE2",X"F6FAFD",X"FBF2F3",X"FFFDFA",X"FCFFFB",X"F2FBFA",X"FBFCFF",X"E8EBF2",X"000505",X"5B6E72",X"EEFDFA",X"FFFCF9",X"FFF9FC",X"FFFBFF",X"F9FFFF",X"FFFAFD",X"FFE6EA",X"D48054",X"D73D01",X"F49569",X"FCFEE9",X"FFFCE9",X"FFF9FA",X"F5FFFF",X"FEF1F8",X"FFFEF8",X"FCFFFF"),
(X"F7F9F6",X"FEFFFF",X"CCE7F8",X"3B75B4",X"295FC1",X"C0DEF8",X"F5FFFA",X"F7FFFF",X"F3F3FB",X"DBE3E5",X"E7F3EF",X"E7F4ED",X"F2F7F1",X"FFFFFD",X"FFFEFF",X"FCFAFD",X"F5FFFF",X"C9DCE2",X"000D0C",X"001402",X"A1D1C3",X"DBFFFF",X"CAFFFF",X"C0FFF6",X"C6FCEF",X"CFF0E9",X"F7FFFF",X"F9FFFD",X"F9FFFF",X"F8FFFF",X"F7FDFD",X"FFFDFF",X"B3F1DC",X"40D4A4",X"097251",X"969F9E",X"FFFDFF",X"FAFAFC",X"FFFBFE",X"FFFEFF",X"FAFDFF",X"FEFDFF",X"FBFAFF",X"FAFFFF",X"FDFEFF",X"FFF8ED",X"F5DA81",X"E2BE10",X"E0AB21",X"D4B855",X"FFF0DE",X"FDF7FF",X"F1FDF1",X"FFFCF6",X"C0AEBE",X"000012",X"727F88",X"FEFCFD",X"E7FFFB",X"CEFFF7",X"AEFFF6",X"9EFFEA",X"D7FFF3",X"F1F4FD",X"FFFFFD",X"FFFDFF",X"F8FFFF",X"F5FFFF",X"E6FFFB",X"88D6C0",X"030D0C",X"555557",X"F8FBFF",X"FFF5FF",X"FCF5FD",X"F5FCFF",X"FFF2FF",X"9C768D",X"000005",X"A9B5B1",X"FBFFFD",X"F6FFF8",X"F0FFF6",X"F8FAF7",X"FFF7FF",X"FFFCFF",X"F7FDFB",X"FFFCFB",X"D9FFED",X"55806C",X"000600",X"EBE9EC",X"FAF7E8",X"D8A458",X"E47E0F",X"FFA23E",X"FFE1E1",X"FFF0F0",X"F3FFFB",X"F2FFFF",X"FDFFFC",X"F8FFFD",X"F5FFFF",X"FFF5FD",X"FEFDFF",X"EDB6D3",X"D9006A",X"C80877",X"FACBEB",X"FFFDFD",X"F1FFFE",X"FBFFFA",X"FFFFF6",X"FCFFF8",X"FBFFF3",X"FBFFEC",X"FDFFF7",X"FFFCFF",X"FDFDFD",X"FAFFE9",X"A7A46F",X"0C0100",X"9B8D9C",X"FBFAFF",X"F5FFFF",X"E0EDFF",X"DBF3FF",X"C4E7FF",X"EBEAF0",X"FDFDFF",X"FBFBFB",X"FDFDFB",X"FFFFFD",X"FCFCFC",X"FFFFFF",X"FEFDFF",X"FFFEFF",X"FEFFFF",X"F9FFFD",X"FFFEFF",X"FFFCFF",X"F9FFFF",X"FFF4F6",X"CE7287",X"AA0001",X"C63552",X"FFD4E7",X"F3FFFF",X"FAFFFC",X"FBFFFF",X"F8FDFF",X"FFFDFA",X"FAFEFD",X"FFFCFF",X"FEF6FF",X"FBFAF8",X"F4FFE7",X"83A96E",X"679E4D",X"56953A",X"D6DFCE",X"F7FFFA",X"FBFFFF",X"F3FCF9",X"F4FFFA",X"DECED1",X"590025",X"A60054",X"FFADDA",X"FFE3FF",X"FFE2FF",X"FFCFEF",X"FFC1EA",X"FFC9EA",X"FEEFF4",X"FFFEFA",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"F8FFFA",X"FFFAFF",X"FFFEFD",X"FDFFF5",X"D4D6E5",X"000825",X"001C2D",X"92A5B4",X"ECFFFF",X"FEFEFF",X"FFF9FD",X"FCFCFC",X"FCFFFF",X"FFFDFF",X"FFFAFE",X"FFFEFB",X"FFFCF9",X"FFFFFD",X"F6FFFC",X"FCFFFB",X"FFECEC",X"9F6E74",X"240006",X"E2D9DA",X"FFFCFD",X"97626C",X"640314",X"923746",X"F5CED1",X"FBFFFB",X"F7FBFA",X"FFF7FE",X"FFFEFA",X"FFF6FF",X"FFF8FF",X"FFEEF5",X"C18086",X"64000C",X"C17E87",X"FCF7F4",X"F6FFFF",X"FEFCFF",X"FFF8FB",X"FFFBFF",X"FEFFFF",X"F8FFFF",X"FFFDFE",X"FFFAFB",X"FFEEFF",X"4A2F40",X"3B2733",X"EBE4EB",X"FFFEFF",X"FDF8FC",X"F9F5F6",X"FCFEFB",X"FBFFFA",X"BEC9E7",X"193684",X"1C59C4",X"0859C4",X"448CDE",X"C2E6FF",X"F9FDFF",X"FAF9FF",X"FFFCFD",X"FFFBFA",X"FFFAFB",X"FFFDFF",X"F9F9F9",X"FCFFFB",X"F8FFF8",X"FAF2FD",X"7C8687",X"080000",X"F8E3E0",X"FFF5FF",X"E38ACC",X"D130A0",X"CF36AA",X"FBDAEB",X"FFFBFF",X"F7FDFD",X"FEFFFF",X"FFFBFC",X"FEFCFD",X"FBFBFD",X"FAFBFD",X"F5B1EC",X"BC1275",X"F0B7DA",X"EAFEF5",X"F0CAEF",X"CB69BE",X"A90983",X"D73CC8",X"F25CCA",X"FFD0FF",X"FEFAFF",X"F4F6F5",X"FAF4F6",X"FFFAFF",X"FFFCFF",X"777E86",X"1B1C55",X"DDE5F8",X"FFFFFB",X"FDFDFB",X"FFFEFF",X"FFFEFF",X"FEFFFF",X"FAEFF7",X"6F6276",X"1D0019",X"E8DAE7",X"FFFAFB",X"DB98CD",X"8C1879",X"E037AE",X"D042B2",X"FFACF7",X"FFEAFF",X"FCFFFF",X"F3F9F7",X"FFFDFB",X"FFFDFB",X"E3E8E2",X"000700",X"7B707E",X"F9FDFE",X"F8FFF8",X"FFFDFC",X"FFF9FF",X"FBFEFF",X"F9FFFD",X"F7F4EF",X"D47F78",X"B41C00",X"FD9067",X"FFF0CF",X"FFEDCA",X"FFDCC5",X"FFD8BC",X"FFE5A2",X"FADACB",X"FFFCEF"),
(X"FEFFFD",X"FDFEFF",X"D0EBFC",X"0E4887",X"073D9F",X"7D9BB5",X"9EA9A3",X"969EAB",X"6A6A72",X"50585A",X"5E6A66",X"CCD9D2",X"FBFFFA",X"FCFCFA",X"F8F6F7",X"FDFBFE",X"F5FFFF",X"DBEEF4",X"5A8685",X"589381",X"97C7B9",X"AFDCD9",X"97D6CE",X"7EC9B4",X"75AB9E",X"88A9A2",X"EFFBF9",X"FBFFFF",X"EDF6F3",X"F2FDF9",X"FBFFFF",X"FFFCFF",X"B3F1DC",X"41D5A5",X"004827",X"959E9D",X"FFFDFF",X"FCFCFE",X"FFF8FB",X"FFFEFF",X"FAFDFF",X"FEFDFF",X"FDFCFF",X"FBFFFF",X"F7F8FD",X"FFF7EC",X"FFEA91",X"E1BD0F",X"EFBA30",X"C4A845",X"FEEDDB",X"FFFCFF",X"F4FFF4",X"FFFEF8",X"C6B4C4",X"020518",X"3B4851",X"9E9C9D",X"82A796",X"83B9AC",X"67C4AF",X"35A881",X"92BCAE",X"FCFFFF",X"FFFFFD",X"FEF8FA",X"F8FFFF",X"F8FFFF",X"E4FDF9",X"78C6B0",X"000302",X"6B6B6D",X"FAFDFF",X"FFE8F7",X"FEF7FF",X"F8FFFF",X"FDDAF0",X"674158",X"5E5F64",X"F2FEFA",X"FBFFFD",X"F6FFF8",X"F3FFF9",X"FBFDFA",X"FFF8FF",X"FFFCFF",X"F4FAF8",X"FFFCFB",X"D2FCE6",X"1A4531",X"8B988E",X"FAF8FB",X"FAF7E8",X"FFD488",X"EC8617",X"CE6804",X"E9C5C5",X"FFFAFA",X"F2FFFA",X"F0FFFD",X"FCFEFB",X"F2FDF7",X"F3FFFD",X"FFFBFF",X"FEFDFF",X"F0B9D6",X"DC006D",X"BF006E",X"FECFEF",X"FFFDFD",X"F0FFFD",X"FBFFFA",X"FEFFF5",X"FCFFF8",X"FBFFF3",X"FBFFEC",X"FCFFF6",X"FFFCFF",X"FEFEFE",X"FCFFEB",X"D0CD98",X"5A4F31",X"524453",X"B1B0B6",X"8F999B",X"828FB1",X"6C84AA",X"3F628C",X"DDDCE2",X"FBFBFD",X"F8F8F8",X"FDFDFB",X"FFFFFD",X"FDFDFD",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FEFFFF",X"F9FFFD",X"FFFDFF",X"FFFAFF",X"F7FFFF",X"FFF4F6",X"CF7388",X"AB0002",X"BB2A47",X"FACFE2",X"F3FFFF",X"FAFFFC",X"FAFEFF",X"F9FEFF",X"FFFDFA",X"FBFFFE",X"FAF7FE",X"FFF9FF",X"FBFAF8",X"F6FFE9",X"ACD297",X"5E9544",X"56953A",X"D3DCCB",X"F4FFF7",X"F7FDFD",X"F2FBF8",X"F4FFFA",X"DDCDD0",X"690835",X"BE186C",X"CD6C99",X"D18BAF",X"AD7091",X"9A5979",X"9C3B64",X"671334",X"EFE0E5",X"FFFFFB",X"FEFEFE",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"F8FFFA",X"FFF5FF",X"FFFEFD",X"FEFFF6",X"D9DBEA",X"1A415E",X"2B6475",X"AFC2D1",X"EEFFFF",X"FFFFFF",X"FFF9FD",X"FCFCFC",X"FCFFFF",X"FFFDFF",X"FFFAFE",X"FFFEFB",X"FFFCF9",X"FCFBF9",X"EDF6F3",X"FCFFFB",X"E5CDCD",X"35040A",X"A27D84",X"FAF1F2",X"FFF8F9",X"DCA7B1",X"5B000B",X"5A000E",X"D7B0B3",X"F7FEF7",X"FCFFFF",X"FFF8FF",X"FFFEFA",X"FFF7FF",X"FFF8FF",X"FFEDF4",X"C28187",X"65010D",X"BA7780",X"F8F3F0",X"F6FFFF",X"FDFBFE",X"FFF8FB",X"FFFAFE",X"FEFFFF",X"F8FFFF",X"FFFDFE",X"FFFAFB",X"FFE6F9",X"44293A",X"422E3A",X"EEE7EE",X"FFFEFF",X"FFFAFE",X"FFFBFC",X"FCFEFB",X"F6FBF5",X"F4FFFF",X"95B2FF",X"0845B0",X"1263CE",X"0D55A7",X"4A6EA0",X"D7DBF8",X"FEFDFF",X"FFFAFB",X"FFFBFA",X"FFFBFC",X"FFFDFF",X"FDFDFD",X"F6FBF5",X"FBFFFB",X"DFD7E2",X"000809",X"9D9290",X"FFF7F4",X"FFF3FF",X"FFAEF0",X"E746B6",X"C42B9F",X"E0BFD0",X"FFFBFF",X"FBFFFF",X"F6F8F7",X"FFFEFF",X"FFFDFE",X"F8F8FA",X"FAFBFD",X"FFBBF6",X"9F0058",X"E0A7CA",X"EFFFFA",X"FFEFFF",X"FFB4FF",X"DB3BB5",X"CB30BC",X"A7117F",X"CD8BC8",X"F7F3FF",X"FEFFFF",X"FFFDFF",X"FEF2FC",X"FFFCFF",X"757C84",X"000033",X"DAE2F5",X"FFFFFB",X"FAFAF8",X"FBFAFF",X"FFFEFF",X"FEFFFF",X"F4E9F1",X"65586C",X"72416E",X"F0E2EF",X"FFF4F5",X"FFD6FF",X"F985E6",X"B40B82",X"ED5FCF",X"9D317C",X"F7C7F1",X"F2F5FE",X"F6FCFA",X"FFFDFB",X"FFF9F7",X"E8EDE7",X"000900",X"7C717F",X"F9FDFE",X"F8FFF8",X"FFFEFD",X"FFFBFF",X"F9FCFF",X"F7FDFB",X"F8F5F0",X"BD6861",X"DC441D",X"E77A51",X"D6BC9B",X"D6AB88",X"D28770",X"B9795D",X"9A611E",X"D0B0A1",X"FFFBEE"),
(X"FBFFFB",X"F3F7F6",X"D9E2DF",X"26322E",X"000600",X"5F696A",X"767F7C",X"7B809E",X"3F4247",X"000204",X"263530",X"EBF8F1",X"F7FDF9",X"FCFEFB",X"FCFCFE",X"FEFFFF",X"FFF9F7",X"C7F2EB",X"50BDA0",X"3ED79E",X"26BA80",X"5DBFA6",X"83CCC5",X"60BCAD",X"27B48A",X"7DDABF",X"EEFFFF",X"FFF5FA",X"FFFAFF",X"FFFEFF",X"F5F6F8",X"F9FFFF",X"B6EFDE",X"5FB298",X"000D0A",X"AA99A1",X"FDFDFD",X"F9FFFF",X"EEFFF9",X"FFFBFF",X"FEFFEC",X"FCFEFD",X"F6FDF5",X"F3FFED",X"F0FEFF",X"FFFCFF",X"FFF3B5",X"CFBF0A",X"F7C526",X"BBAA28",X"F8E9D2",X"FFFDFF",X"F5FFF2",X"FDFCFF",X"D0AACF",X"2E0044",X"63426D",X"6E6C71",X"6F8171",X"86C1AD",X"55C1A9",X"2AAC8A",X"7DE1C5",X"E2FFFF",X"FFF8FB",X"FFF5F9",X"FFFDFF",X"FFFBFF",X"E9FFFF",X"7EC9B5",X"000106",X"485254",X"FFCBFF",X"FFC4FF",X"FFB6FF",X"FF99FF",X"F455C9",X"BE62AD",X"E6D8EF",X"FFFCFD",X"FBFFF1",X"FAFDF2",X"F6FFF8",X"FCFBFF",X"FFF7FF",X"FAFDFF",X"ECFFFC",X"FDFFF9",X"B1E5BF",X"0D2611",X"D5D1CE",X"FFF6FC",X"FFF7E9",X"FFE1A0",X"E5A34C",X"A56122",X"687269",X"FFFFFD",X"F8FCFB",X"FBFAF8",X"FFF9FA",X"FFFBF8",X"F9FDFE",X"FFF8FF",X"FFFAFF",X"FFB5E1",X"D60266",X"8C093D",X"F0DBD8",X"FFF6FF",X"F2FDFF",X"FFFCFF",X"FFFBFF",X"FFFCFF",X"FFFEFF",X"FEFEF4",X"FFFCF3",X"FFFBFF",X"FFFBFE",X"FFFCF2",X"E5D452",X"C9B022",X"220800",X"000000",X"698289",X"5B7C9F",X"0D4381",X"2675D1",X"E7E6EC",X"FFFEFF",X"FAFAFC",X"FCFCFA",X"FFFFFD",X"FCFCFA",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"FAFFFC",X"FDFFFE",X"FFFAFE",X"FAFEFF",X"FFF2F5",X"CD7486",X"9D0105",X"CB123B",X"FFC0D9",X"FAFEFF",X"FEFFFF",X"F3FFFF",X"FEFFFF",X"FFFDFD",X"FBFFF8",X"FBFBF3",X"FFFCFB",X"FFFBFA",X"F5FDF0",X"C8E8C1",X"5E964F",X"509538",X"CDDECB",X"F2FFF6",X"FDFBFC",X"FAFAFA",X"F9FFFD",X"F9BFD7",X"980148",X"CC1572",X"B85486",X"B37398",X"AF80A4",X"B26A9C",X"A00956",X"A5054F",X"FFD8EE",X"EAFFF6",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FBFFF9",X"F8FAF9",X"F0FFFD",X"F5FFFF",X"CEF7FF",X"0894C9",X"04A7E0",X"7FC7F7",X"EEFFFF",X"FFFEFF",X"FFF9F9",X"FCFDF8",X"FBFFFF",X"FFFEFF",X"FEFCFF",X"FBFFFF",X"F5FFF6",X"F5FAF3",X"FFFCFB",X"FFEAEF",X"E29EA9",X"53000B",X"EAA4AF",X"FFF0F2",X"FFF2F0",X"FFDFE2",X"953843",X"740012",X"A95263",X"FFE8ED",X"F5F1EE",X"FFFCF9",X"EEFFFD",X"FFFEFF",X"FCFBFF",X"F7F9F6",X"AB8884",X"5F0912",X"AF6973",X"FFF1F0",X"FFFCFF",X"FFFAFE",X"FFFBFB",X"FFFCFE",X"FFFDFF",X"FDFEFF",X"F6FFFE",X"F2FFFB",X"F1ECF0",X"282A36",X"3B3E51",X"EAE7F8",X"FDFCFF",X"FBFFFA",X"FFFFFD",X"FFFAFF",X"F8FDFF",X"F9FCF1",X"F4FCEF",X"9CB7CC",X"00337F",X"1D67D4",X"0457BF",X"2579CF",X"C0F3FF",X"EBFFFF",X"F9FAF2",X"FFFFFF",X"FFFBFC",X"FFF5F2",X"FFFCF9",X"F4FFFF",X"B7BAE3",X"000013",X"A38F9A",X"FFFAFF",X"EEFEFD",X"D6C8D5",X"7F4168",X"6A3263",X"897689",X"FFF5FF",X"FFFBFF",X"FAFCF7",X"FFFFFA",X"FFF8F9",X"FFFFFF",X"F2FFFF",X"DAC1D7",X"0B0010",X"9AA698",X"FFFFEF",X"F6F8F7",X"F9FDFF",X"F7C7E1",X"AA438A",X"D42BBA",X"B7088B",X"F778D3",X"FFE4FF",X"FCFBF9",X"F4F6F1",X"FFF6FF",X"B89BB9",X"330028",X"F1E3F4",X"FFFEF8",X"FBFDFC",X"FDFBFF",X"FFFCFF",X"F8FFFF",X"FFDEF1",X"C163B9",X"B10077",X"FFD4FF",X"FFFCFD",X"F5F7F4",X"FFEFFF",X"BD7EAB",X"A01D7A",X"E12F9D",X"760F56",X"E6CEE8",X"F7FFFF",X"EEFFFB",X"F2FFF8",X"EEEEEC",X"0A0000",X"7E717B",X"F9FDFE",X"F7FFFC",X"FFFFFD",X"FFFEFF",X"F9FEFF",X"F7FFFE",X"FAFCF7",X"636B6E",X"7B502E",X"AE7655",X"C19C8A",X"C4A589",X"C0997C",X"C67B5C",X"C54A0F",X"D3A595",X"FFF9EA"),
(X"EFF6EF",X"FCFFFF",X"DFE8E5",X"3D4945",X"000600",X"C5CFD0",X"F9FFFF",X"F5FAFF",X"ECEFF4",X"C2CACC",X"52615C",X"D5E2DB",X"FBFFFD",X"F6F8F5",X"FFFFFF",X"F4F5F7",X"FFFCFA",X"C8F3EC",X"00674A",X"008F56",X"52E6AC",X"A8FFF1",X"C5FFFF",X"AAFFF7",X"55E2B8",X"7AD7BC",X"E1FAF4",X"FFF9FE",X"FFF6FB",X"FFFCFD",X"FEFFFF",X"F8FEFE",X"B4EDDC",X"42957B",X"000502",X"AF9EA6",X"FCFCFC",X"F9FFFF",X"EFFFFA",X"FFFBFF",X"FDFFEB",X"FBFDFC",X"FAFFF9",X"F4FFEE",X"F3FFFF",X"FEFBFF",X"FFF2B4",X"D4C40F",X"F0BE1F",X"C4B331",X"F6E7D0",X"FFFAFC",X"F3FFF0",X"F9F8FF",X"CAA4C9",X"3A0450",X"94739E",X"FDFBFF",X"F2FFF4",X"D1FFF8",X"9DFFF1",X"5DDFBD",X"7ADEC2",X"DFFFFE",X"FFF5F8",X"FFFAFE",X"FFFDFF",X"FDF3FB",X"ECFFFF",X"8BD6C2",X"0D0E13",X"000709",X"733A6F",X"B359A1",X"89217A",X"C941AF",X"E041B5",X"EC90DB",X"FFF6FF",X"FFF7F8",X"FAFEF0",X"FCFFF4",X"F5FFF7",X"FDFCFF",X"FFF4FF",X"FAFDFF",X"F1FFFF",X"F3F6EF",X"95C9A3",X"334C37",X"8C8885",X"BFACB2",X"E7CABC",X"EDBA79",X"E3A14A",X"813D00",X"010B02",X"D4D4D2",X"FBFFFE",X"FFFFFD",X"FFFAFB",X"FFFEFB",X"F9FDFE",X"FFF5FF",X"FFFAFF",X"FFB4E0",X"CE005E",X"780029",X"EFDAD7",X"FFF6FF",X"F4FFFF",X"FFFCFF",X"FFFBFF",X"FFFBFF",X"FFFDFF",X"FDFDF3",X"FFFCF3",X"FFFCFF",X"FFFAFD",X"FFFBF1",X"DBCA48",X"D8BF31",X"9D8348",X"DBDBD9",X"E5FEFF",X"D2F3FF",X"9CD2FF",X"2271CD",X"EDECF2",X"FFFEFF",X"FDFDFF",X"FEFEFC",X"FFFFFD",X"FDFDFB",X"FFFFFF",X"FFFFFF",X"FFFEFF",X"FFFDFE",X"FAFFFC",X"FDFFFE",X"FFFCFF",X"FCFFFF",X"FFF3F6",X"CD7486",X"9E0206",X"C10831",X"FFBCD5",X"FAFEFF",X"FEFFFF",X"F3FFFF",X"FEFFFF",X"FFFDFD",X"FBFFF8",X"FFFFF7",X"FFFAF9",X"FFFAF9",X"FBFFF6",X"BBDBB4",X"639B54",X"498E31",X"CFE0CD",X"F4FFF8",X"FFFEFF",X"FCFCFC",X"F9FFFD",X"F7BDD5",X"9A034A",X"B7005D",X"FFAFE1",X"FFD8FD",X"FFE3FF",X"FFD1FF",X"FF91DE",X"9F0049",X"FFD5EB",X"F1FFFD",X"FDFDFD",X"FDFDFD",X"FEFEFE",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FAFFF8",X"FEFFFF",X"EFFFFC",X"F0FFFA",X"CEF7FF",X"0D99CE",X"009DD6",X"73BBEB",X"ECFFFE",X"FFFEFF",X"FFFAFA",X"FCFDF8",X"FBFFFF",X"FFFEFF",X"FDFBFF",X"FBFFFF",X"F2FFF3",X"FCFFFA",X"FDF3F2",X"FFE5EA",X"712D38",X"620A1A",X"BF7984",X"D0ACAE",X"CDB5B3",X"B88689",X"7B1E29",X"881326",X"5C0516",X"E7C7CC",X"FFFEFB",X"FFFEFB",X"F0FFFF",X"FFFEFF",X"FBFAFF",X"F9FBF8",X"A78480",X"57010A",X"914B55",X"FBEDEC",X"FFFCFF",X"FFFBFF",X"FFFBFB",X"FFFDFF",X"FFFDFF",X"FDFEFF",X"F6FFFE",X"F2FFFB",X"F2EDF1",X"191B27",X"424558",X"EBE8F9",X"FFFEFF",X"FBFFFA",X"FFFFFD",X"FFFBFF",X"FBFFFF",X"FBFEF3",X"FBFFF6",X"E8FFFF",X"89BEFF",X"0953C0",X"1E71D9",X"0155AB",X"5C8FA0",X"E6FBFC",X"FFFFF8",X"F8F8F8",X"FFFDFE",X"FFF6F3",X"FFFEFB",X"E8F5FE",X"6E719A",X"000519",X"55414C",X"A0939A",X"899998",X"362835",X"2B0014",X"2E0027",X"0E000E",X"E8DAE7",X"FFFBFF",X"F9FBF6",X"FEFDF8",X"FFF7F8",X"FDFDFF",X"F5FFFF",X"D6BDD3",X"0D0212",X"A4B0A2",X"FDFFED",X"F8FAF9",X"FCFFFF",X"FFEAFF",X"FFA6ED",X"AC0392",X"F344C7",X"9E1F7A",X"CD9EC2",X"FCFBF9",X"F7F9F4",X"FFFAFF",X"D6B9D7",X"601055",X"F6E8F9",X"FFFDF7",X"FDFFFE",X"FFFDFF",X"FEF7FF",X"F7FFFF",X"FFE1F4",X"C668BE",X"C20988",X"F6C6FA",X"FCF3F4",X"FDFFFC",X"FFEEFE",X"FFDFFF",X"EE6BC8",X"B80674",X"5D003D",X"100012",X"C9D5D5",X"EEFFFB",X"F7FFFD",X"EFEFED",X"0D0001",X"7E717B",X"FAFEFF",X"F7FFFC",X"FFFFFD",X"FDFBFE",X"F9FEFF",X"F8FFFF",X"FDFFFA",X"6B7376",X"220000",X"CC9473",X"FFF6E4",X"FFE3C7",X"FFEACD",X"FFD2B3",X"F0753A",X"DCAE9E",X"FFF8E9"),
(X"FFFFF4",X"F7FBE2",X"FAF7D8",X"BBB257",X"989A00",X"DCDEAC",X"FCFEFB",X"F3EFF0",X"FCFBFF",X"FBFFFF",X"CCD7D3",X"E9F2ED",X"F9FEFA",X"FDFDFD",X"FEFEFF",X"FEFFFF",X"FFF9F2",X"D1E3EF",X"00031B",X"000207",X"B8C3B3",X"FFFFF6",X"FEF5FA",X"F0FFFF",X"DFFEF9",X"D1ECE7",X"F2F6F7",X"FFFCFF",X"FBFFFF",X"F4FFFB",X"F7FDFD",X"F3FFFF",X"B7E5DA",X"3B6156",X"000002",X"A3A3A3",X"FDFFFE",X"FFFDFE",X"FCFDFF",X"FFF8FF",X"FFF8FF",X"FFF6FF",X"FFFBFF",X"FFFFF2",X"FFFEFB",X"FFF3F5",X"FFE591",X"E6C000",X"E0C216",X"D4CE76",X"FEF7ED",X"FFFEF5",X"F8FFFF",X"FEF4FF",X"D895D8",X"69006C",X"8E529A",X"F1F7FF",X"FBFBEF",X"FCFEF9",X"F7F9FF",X"D9DDE6",X"C3E4DD",X"FFFAFF",X"EEFFFB",X"FEFFFF",X"FBFFFF",X"FEF3FB",X"E6FFFF",X"91D5C6",X"003A2C",X"030009",X"B69BAA",X"EFCBE7",X"C887C1",X"BF49A9",X"EE4BC0",X"F659C2",X"FFBFFA",X"FFF7FF",X"FFF6FF",X"FFFEFF",X"FDF7F9",X"FFFCFF",X"FCF9FF",X"FFF8FF",X"F5FFFF",X"AEEFD9",X"7AB285",X"394434",X"080000",X"250908",X"CF997F",X"D3A16C",X"5E4E2A",X"0B0813",X"03000B",X"BF9DB5",X"FFF6FF",X"FDFEFF",X"FEFAF9",X"FFFCFB",X"FFFDFE",X"FFFCFF",X"FFFCFA",X"FCADCC",X"8D073A",X"28030A",X"D4E8CF",X"FFF9F3",X"FFFEF9",X"FFFFF3",X"FEFFE5",X"FFFEFC",X"FEF9FF",X"FDFBFF",X"FCFCFF",X"FFFEFF",X"FFFDF8",X"FFFBE5",X"E5C95B",X"D5B009",X"EBC66B",X"F9F0EB",X"FBFFFD",X"FFFDF6",X"FBFFFD",X"B3D5DE",X"F1F0F8",X"F9F8FE",X"FDFDFF",X"FFFFFF",X"FFFFFD",X"FFFFFD",X"FEFEFC",X"FCFCFC",X"FFFEFF",X"FFFDFE",X"F9FFFB",X"FBFFFF",X"FFFDFF",X"FFFFFF",X"FFF1F4",X"C57483",X"9E0605",X"BE0121",X"FEBFC8",X"FFFCF9",X"FFF6FF",X"F7FFFF",X"FFFDFF",X"FFFAFF",X"FAFFF8",X"FFFFFB",X"FFFBFC",X"F8FAF7",X"F5FFF6",X"98BB9A",X"609261",X"5D975C",X"D8E3D5",X"F4FEF6",X"FFF2FB",X"FFF6FF",X"FDFEFF",X"FFB4DD",X"AD0359",X"A70261",X"F5A4CF",X"FFF3FF",X"FAF4FF",X"F3F3FF",X"FFF9FF",X"C099B6",X"F8E6F2",X"FCFFFB",X"FDFDFD",X"FDFDFD",X"FEFEFE",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFF4FA",X"FFF7FF",X"FFF9FF",X"FFFAFF",X"C9ECFF",X"009AE4",X"00A3F9",X"7BBDFA",X"E6FEFF",X"FDFDFF",X"FFFBFD",X"FFFCF6",X"FFFFF6",X"FFFCF3",X"FFFAF1",X"FFFFF1",X"FFFAFB",X"F7F7F7",X"FFFFFF",X"D2BBC3",X"391119",X"351113",X"1A0000",X"2B060D",X"390511",X"866C6B",X"826662",X"480F16",X"480A19",X"A48A93",X"FEFFFF",X"F4F5F7",X"FFFDFF",X"F4FFFF",X"EFFFFF",X"FBFBF9",X"9C8786",X"1D0302",X"4A3C3C",X"EDECF1",X"FFFAFF",X"FCFDFF",X"F5FFFB",X"F9FFFF",X"FFFDFF",X"FFFAFF",X"FAFEFF",X"F4FFFD",X"D1D2CD",X"00030C",X"404C64",X"E7E5FD",X"FEFDFF",X"F6FFF6",X"FCFFFB",X"FFFAFF",X"FDFCFA",X"FFFFFD",X"F8F9F4",X"FAFCF9",X"EEF6FF",X"8BA7CF",X"1D529E",X"266ED4",X"0546A4",X"99BFFF",X"F4FFFF",X"F4F2FF",X"FFFCFF",X"FFFBFF",X"FBFCFF",X"C2D2F4",X"26478E",X"00092B",X"373E46",X"444245",X"0A150F",X"010800",X"00040B",X"00394C",X"000D1B",X"8E9FAF",X"FCF9FF",X"F8F8F6",X"FCFDF7",X"FFFAF8",X"FBF6FA",X"F7FFFF",X"DBBCDE",X"000023",X"B5A4C6",X"FFF2FF",X"FFF9FF",X"FFFEFF",X"FBF8EF",X"FFF0F8",X"EABDDE",X"9E247B",X"DB2BB2",X"AD0089",X"FF93FD",X"FFE1FF",X"FEF3FF",X"EBCFDB",X"A41072",X"FFDBFA",X"FFF9F9",X"FBFFFC",X"FFFEFF",X"FFF6FC",X"F7FFFF",X"FFD7FB",X"C82797",X"CC0288",X"FCCDFF",X"FFF9FF",X"EFFFFF",X"F1F7F3",X"FFF7FF",X"FFD5FF",X"926085",X"2C001C",X"251021",X"222F35",X"C2DADE",X"F7FEFF",X"F2EFFA",X"000005",X"717777",X"F7FFFD",X"FCFEFB",X"FFFBFD",X"F9FAFC",X"F5FFFF",X"FFFEFF",X"FFF1FA",X"6C5A66",X"060A00",X"7B7C6C",X"FAE7ED",X"FFFDFB",X"F8FFFF",X"FFFFFD",X"EACAB5",X"E8CDC4",X"FFF9F3"),
(X"FFFDF2",X"FEFFE9",X"F7F4D5",X"E9E085",X"E8EA49",X"ECEEBC",X"FAFCF9",X"FFFDFE",X"FFFEFF",X"EDF3F3",X"F8FFFF",X"F5FEF9",X"FAFFFB",X"FDFDFD",X"FCFCFE",X"FAFBFD",X"FFFDF6",X"C7D9E5",X"071931",X"000308",X"BAC5B5",X"FFFFF6",X"FCF3F8",X"E8FDFE",X"E4FFFE",X"EDFFFF",X"FCFFFF",X"FFF7FA",X"F8FEFC",X"F8FFFF",X"F8FEFE",X"EFFFFC",X"B4E2D7",X"22483D",X"030406",X"A1A1A1",X"FEFFFF",X"FBF9FA",X"FEFFFF",X"FFF7FF",X"FFFBFF",X"FFF5FF",X"FFF9FF",X"FCFAED",X"FFFEFB",X"FFF5F7",X"FDDA86",X"DBB500",X"DABC10",X"E9E38B",X"FFFEF4",X"FFFCF3",X"F5FFFE",X"FAF0FF",X"CF8CCF",X"68006B",X"7D4189",X"E1E7F3",X"FBFBEF",X"FEFFFB",X"F7F9FF",X"FBFFFF",X"E9FFFF",X"FFF2F9",X"F0FFFD",X"FBFDFC",X"F9FFFF",X"FFFAFF",X"E3FFFC",X"8BCFC0",X"0D5547",X"3D3743",X"F9DEED",X"FFE7FF",X"FFDEFF",X"FF90F0",X"D532A7",X"DE41AA",X"C974AF",X"F2E3F6",X"FFF3FD",X"FFFEFF",X"FAF4F6",X"FFFCFF",X"FCF9FF",X"FEF6FF",X"EFFDFD",X"92D3BD",X"74AC7F",X"8E9989",X"D9CDCF",X"EED2D1",X"FFE7CD",X"FFEBB6",X"DBCBA7",X"191621",X"03000B",X"87657D",X"F9E2F4",X"FBFCFF",X"FFFCFB",X"FFFAF9",X"FFFDFE",X"FEFBFF",X"FFFCFA",X"F5A6C5",X"80002D",X"1C0000",X"D4E8CF",X"FFF7F1",X"FDFCF7",X"FFFFF3",X"FFFFE6",X"FFFFFD",X"FEF9FF",X"FDFBFF",X"FDFDFF",X"FFFEFF",X"FFFDF8",X"FFFAE4",X"D9BD4F",X"D6B10A",X"F7D277",X"FFFBF6",X"F7FDF9",X"FCF9F2",X"F1F7F3",X"E6FFFF",X"FFFEFF",X"FBFAFF",X"FEFEFF",X"FEFEFE",X"FCFCFA",X"FFFFFD",X"FFFFFD",X"FFFFFF",X"FFFEFF",X"FFFEFF",X"F9FFFB",X"FBFFFF",X"FFFDFF",X"FEFEFE",X"FFEEF1",X"C06F7E",X"A00807",X"BB001E",X"FDBEC7",X"FFFCF9",X"FFF6FF",X"F7FFFF",X"FFFDFF",X"FFF9FE",X"F9FEF7",X"FFFFFB",X"FFFEFF",X"F6F8F5",X"F2FFF3",X"84A786",X"588A59",X"7DB77C",X"F1FCEE",X"F9FFFB",X"FFF1FA",X"FFFAFF",X"FDFEFF",X"FEADD6",X"AC0258",X"A80362",X"EC9BC6",X"FFF0FF",X"FFFCFF",X"FCFCFF",X"F8ECFF",X"FFF0FF",X"FFF8FF",X"F8FDF7",X"FDFDFD",X"FDFDFD",X"FDFDFD",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FFF8FE",X"FFF1F9",X"FFF8FF",X"FFFBFF",X"C1E4FF",X"019DE7",X"00A7FD",X"64A6E3",X"E4FCFF",X"FCFCFF",X"FFFBFD",X"FFFDF7",X"FFFFF6",X"FFFCF3",X"FFF9F0",X"FFFFF1",X"FFF5F6",X"FCFCFC",X"FDFDFF",X"836C74",X"1B0000",X"795557",X"E5C5C6",X"F5D0D7",X"FFD5E1",X"FFEFEE",X"FFE9E5",X"8F565D",X"2A0000",X"442A33",X"E4E5E9",X"FEFFFF",X"FFFCFF",X"EDFBFC",X"F1FFFF",X"FCFCFA",X"A08B8A",X"120000",X"392B2B",X"F1F0F5",X"FFFAFF",X"FDFEFF",X"F6FFFC",X"F9FFFF",X"FFFDFF",X"FFFAFF",X"FAFEFF",X"F3FFFC",X"C3C4BF",X"00030C",X"57637B",X"F0EEFF",X"FFFEFF",X"F7FFF7",X"FBFFFA",X"FFF8FF",X"FFFEFC",X"FDFDFB",X"FFFFFB",X"FEFFFD",X"F8FFFF",X"DCF8FF",X"4F84D0",X"0C54BA",X"1B5CBA",X"4369AA",X"E4EFFF",X"FFFDFF",X"FCF5FC",X"FFF9FF",X"F5F6FF",X"9FAFD1",X"000F56",X"91AFD1",X"DDE4EC",X"F2F0F3",X"E0EBE5",X"CED5CD",X"B1C0C7",X"5A93A6",X"4D7E8C",X"3E4F5F",X"F0EDF8",X"FFFFFD",X"FBFCF6",X"FFF9F7",X"FFFDFF",X"F6FFFF",X"D8B9DB",X"090830",X"B8A7C9",X"FFF5FF",X"FFF7FF",X"F5F3F8",X"FFFFF6",X"FFEAF2",X"FFEBFF",X"FF9EF5",X"D424AB",X"D825B4",X"9B127C",X"E3ABDC",X"FFFAFF",X"E4C8D4",X"A10D6F",X"FCD7F6",X"FFFBFB",X"FBFFFC",X"FFFEFF",X"FFF8FE",X"F7FFFF",X"FFD0F4",X"DA39A9",X"C90085",X"FCCDFF",X"FFF1FE",X"F0FFFF",X"FBFFFD",X"FFF2FF",X"FFE9FF",X"FFCFF4",X"4F223F",X"0D0009",X"0A171D",X"3A5256",X"E5ECF6",X"EEEBF6",X"010207",X"717777",X"F8FFFE",X"FDFFFC",X"FFFCFE",X"FCFDFF",X"F7FFFF",X"FFFDFE",X"FFEBF4",X"715F6B",X"000400",X"5F6050",X"FBE8EE",X"FFFDFB",X"F2FDF9",X"F9F8F6",X"FFF6E1",X"FFF7EE",X"FFFCF6"),
(X"FFFAFE",X"FFFEFF",X"FBEDD3",X"FEE45C",X"E7D904",X"EDE4A3",X"FFFEFF",X"FFF9F7",X"FFFAFE",X"FCFCFC",X"FCFEFD",X"FCFEFD",X"FEFCFD",X"FFFCFD",X"FDFBFE",X"FCFCFE",X"FFFEFD",X"B3E4FF",X"3765A1",X"00002C",X"BEC3C6",X"FCFFF1",X"FBF8F1",X"FEFFFF",X"FFF5FF",X"F5FFFF",X"F5FEFD",X"FFFCFE",X"FFFDFF",X"FFF4FA",X"FFF6FE",X"EFFEFB",X"AED9CF",X"242529",X"040507",X"9C9E9D",X"FCFAFD",X"FAFFFF",X"FFFEFF",X"F6FEFF",X"F5FFFF",X"F1FBFD",X"FCFFFF",X"FAFDF4",X"FFFEF1",X"FFFED9",X"E8CB67",X"E4BD1A",X"D9B962",X"F3E7DB",X"FFFCFF",X"FBF5F5",X"F8FFFF",X"FEF5FF",X"C67BCD",X"760070",X"7A1C7A",X"EBD2F2",X"F5FFFA",X"FCFCFA",X"FFF3FF",X"FBFEFF",X"F6FFF9",X"FEFBF6",X"FEFFFF",X"FFF6FF",X"FFFFFF",X"FFFFFF",X"CFFFF8",X"49DCB2",X"12BC8D",X"3F6E68",X"EDF9ED",X"F7FFF6",X"F1FDF3",X"F8EBF5",X"EFAFE1",X"B8469E",X"D149B8",X"FF7CF4",X"FFDAFF",X"FBF1FF",X"EEFFFF",X"F5FFFB",X"FEFDFB",X"FAF9FE",X"C4FFFB",X"33DFAF",X"47A581",X"DEFAE4",X"FDFEF6",X"F9FEF8",X"FFFEF4",X"FFFCF0",X"FEFFFF",X"A088A2",X"860044",X"A50054",X"FFA6E5",X"FFF2FF",X"F6FFFF",X"FFFCFD",X"FFF8F9",X"F9FFFF",X"FBFEF3",X"CDA9AD",X"230511",X"000010",X"DBE8F9",X"FCFBFF",X"FFFFFF",X"F4FDFF",X"FCFFFF",X"FAFAFF",X"FBFCFE",X"FBFFFA",X"F7FFFC",X"F7FFFF",X"FCFFF4",X"F7F9D2",X"E4C72E",X"E0BC06",X"E6C96D",X"FBFEED",X"F6FFFA",X"FFF4FE",X"FFF7FF",X"FBFFFF",X"FDFCFF",X"F6F5FA",X"FBFBFD",X"FFFFFF",X"F7F7F7",X"FFFFFD",X"FFFFFD",X"FFFFFD",X"FDFCFF",X"FFFCFE",X"FBFFFC",X"F9FFFD",X"FDFBFC",X"FFFEFF",X"FCE9EB",X"AF717C",X"A90307",X"BA000F",X"F4C5BB",X"F5FFF8",X"FFF5FB",X"FFFFFD",X"FFF7F8",X"FFFDFF",X"FFFEFF",X"FDFDFF",X"F3FCFF",X"F1FFF6",X"CFF5C4",X"73A161",X"5B834E",X"99BC94",X"FCF8F7",X"FFFFFF",X"FFF6FF",X"FDFDFF",X"F1F9FF",X"F39CD1",X"B3015F",X"AC0869",X"E287B3",X"FFF0F9",X"FFF6ED",X"FFFFF3",X"F4FEF6",X"FDFEFF",X"FCFAFF",X"FFF5FE",X"FFFFFF",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"F5FEFF",X"FFF9FF",X"FDFAFF",X"F8FFFF",X"B3EFFA",X"029ED9",X"009CE3",X"5AACD1",X"E4FBFF",X"F8FBFF",X"FFFDFE",X"F9FFFF",X"F1FFFF",X"F7FFFF",X"F9FFFF",X"F0FDFF",X"F9FEFF",X"FDFBFF",X"E0C8E0",X"1B000B",X"160006",X"D6D2D3",X"F7FDFB",X"FFFEFF",X"FFFEFF",X"FCFBF9",X"FFF9F8",X"9E808A",X"24000B",X"22000C",X"C19FBA",X"FFF5FF",X"F9FDFF",X"FFFEFF",X"F9F7FA",X"FFFFFF",X"B197A0",X"260007",X"2A0013",X"E4C3E2",X"FDFDFF",X"F8F9FD",X"FCFFFF",X"F6FFFE",X"F9FFFF",X"FFFEFF",X"FFF4FB",X"FFF6FD",X"AAA5A2",X"00020B",X"5E667D",X"FAF6FF",X"FAF8FD",X"F8FFF8",X"F8FFFA",X"FFF6FF",X"F5FFFF",X"F4FBFF",X"FFFCFF",X"FEEFF6",X"FFFBF4",X"FCFEFD",X"C0DFFB",X"1F568C",X"246CB8",X"18538F",X"D3F2FF",X"FCFFFB",X"FEFFEF",X"EEFDF8",X"D7F0F5",X"334C53",X"464F78",X"DBE9F4",X"FBFFFD",X"FFFEFF",X"FBFAFF",X"FFFBFF",X"EAFCFF",X"93D2E4",X"30B0B3",X"003B4A",X"B1B8CA",X"FFFCFF",X"F7F9F4",X"FFFEFA",X"FFFAFD",X"FCF7FD",X"D3A9E8",X"861986",X"CF96DA",X"F9F8FD",X"FFFBFF",X"FAF8FF",X"F5FEFF",X"FDFBFF",X"EAFFEF",X"FFF6FF",X"F0B3EC",X"9E1E8B",X"DB21B0",X"A5027F",X"FFABFA",X"FFBCEE",X"B40882",X"FFD1FF",X"FFFBFF",X"FBFFF8",X"FFFFFA",X"FFFDFB",X"F6FFFF",X"FFC8F9",X"E116B0",X"C40590",X"FFCDFF",X"FFFCFF",X"FFF8FF",X"FEFFFD",X"FFFAF4",X"F8FBFF",X"FFFDF6",X"D2CFCA",X"000A08",X"053736",X"03363A",X"647C86",X"D2D5DA",X"010000",X"78706E",X"FEFEFC",X"F9F7F8",X"FFF9FC",X"FFFEFF",X"F7FDFB",X"FFFCFF",X"FFE6F4",X"705252",X"050500",X"43464F",X"E5DDEC",X"FFFDFF",X"FFF9FF",X"F8F2FF",X"FAFFFF",X"FFFFF8",X"FEFAF7"),
(X"FFF9FD",X"FFFEFF",X"F7E9CF",X"EAD048",X"EBDD08",X"F0E7A6",X"FFFEFF",X"FEF6F4",X"FFFAFE",X"FDFDFD",X"FCFEFD",X"FDFFFE",X"FFFDFE",X"FFFDFE",X"FEFCFF",X"FDFDFF",X"FAF6F5",X"B3E4FF",X"4775B1",X"000332",X"BABFC2",X"FBFFF0",X"FFFEF7",X"F9FAFC",X"FFF8FF",X"EFFDFD",X"F9FFFF",X"FBF5F7",X"FFFDFF",X"FFF9FF",X"FFF9FF",X"F3FFFF",X"97C2B8",X"040509",X"000002",X"9EA09F",X"FFFEFF",X"F8FEFE",X"FBFAFF",X"F9FFFF",X"F5FFFF",X"F8FFFF",X"FCFFFF",X"FBFEF5",X"FFFEF1",X"FFF4CF",X"ECCF6B",X"ECC522",X"EACA73",X"FFFDF1",X"FDF6FE",X"FDF7F7",X"F8FFFF",X"F5ECFF",X"C075C7",X"7C0376",X"5D005D",X"E7CEEE",X"F0FFF5",X"FDFDFB",X"FFF9FF",X"F0F3F8",X"F3FEF6",X"FFFFFA",X"FBFDFC",X"FFEFF8",X"FAFAFC",X"FAFAFC",X"C5FBEE",X"53E6BC",X"1EC899",X"7BAAA4",X"EEFAEE",X"F7FFF6",X"F8FFFA",X"FFFAFF",X"FFD9FF",X"F785DD",X"CC44B3",X"D64FC7",X"E4A9DF",X"FFF6FF",X"F2FFFF",X"F3FFF9",X"FCFBF9",X"EFEEF3",X"A5ECDC",X"08B484",X"7FDDB9",X"E6FFEC",X"FAFBF3",X"FAFFF9",X"FFFDF3",X"FEFAEE",X"FEFFFF",X"ECD4EE",X"960554",X"B81067",X"CF61A0",X"FFF6FF",X"F6FFFF",X"FFF5F6",X"FFFCFD",X"F4FDFA",X"F9FCF1",X"B18D91",X"1A0008",X"000212",X"C9D6E7",X"FFFEFF",X"F7F7F7",X"F8FFFF",X"F8FBFF",X"FCFCFF",X"FEFFFF",X"F1F8F0",X"F8FFFD",X"F8FFFF",X"F3F9EB",X"F3F5CE",X"E0C32A",X"DEBA04",X"ECCF73",X"FCFFEE",X"F5FFF9",X"FFFAFF",X"FFF6FF",X"F5F9FA",X"FDFCFF",X"FFFEFF",X"FFFFFF",X"F8F8F8",X"FFFFFF",X"FFFFFD",X"F9F9F7",X"FFFFFD",X"FFFEFF",X"FFFCFE",X"FAFFFB",X"F8FFFC",X"FEFCFD",X"FFFEFF",X"FFF1F3",X"91535E",X"AB0509",X"B8000D",X"E6B7AD",X"F3FFF6",X"FFF8FE",X"F9F8F6",X"FFFCFD",X"FFFDFF",X"FBFAFF",X"FBFBFF",X"F8FFFF",X"E9FFEE",X"A5CB9A",X"5B8949",X"769E69",X"CFF2CA",X"FFFEFD",X"FBFBFB",X"FFF4FE",X"FEFEFF",X"F3FBFF",X"E38CC1",X"AC0058",X"AD096A",X"DF84B0",X"FFF4FD",X"FEF5EC",X"FFFCF0",X"F4FEF6",X"FAFBFF",X"FFFEFF",X"FFF1FA",X"FEFEFE",X"FDFDFD",X"FDFDFD",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"F8FFFF",X"FFFCFF",X"F7F4FB",X"F0FBF7",X"ADE9F4",X"029ED9",X"00A5EC",X"4698BD",X"E0F7FD",X"FBFEFF",X"FFFBFC",X"ECF5F2",X"F4FFFF",X"F8FFFF",X"F2F9FF",X"F5FFFF",X"F7FCFF",X"FDFBFF",X"B9A1B9",X"2F041F",X"8A697A",X"F6F2F3",X"F9FFFD",X"FFFDFF",X"FFFEFF",X"F9F8F6",X"FFF9F8",X"EDCFD9",X"35031C",X"471131",X"704E69",X"F6E9FD",X"FAFEFF",X"FCFAFF",X"FFFEFF",X"FBFBFB",X"C4AAB3",X"420A23",X"400929",X"B190AF",X"FDFDFF",X"FAFBFF",X"F6FAF9",X"F9FFFF",X"F3FBFD",X"F4F3F9",X"FFFAFF",X"FFF3FA",X"A7A29F",X"00020B",X"929AB1",X"FBF7FF",X"FFFEFF",X"F5FFF5",X"F6FFF8",X"FFFAFF",X"C7D4DC",X"E3EAFC",X"FBF8FF",X"FFFAFF",X"FEEFE8",X"FBFDFC",X"E6FFFF",X"659CD2",X"003A86",X"124D89",X"D0EFFF",X"FBFFFA",X"FDFEEE",X"F5FFFF",X"99B2B7",X"00070E",X"7881AA",X"F4FFFF",X"F7FDF9",X"F6F5FA",X"FFFEFF",X"FFFDFF",X"EBFDFF",X"ADECFE",X"38B8BB",X"1B5A69",X"545B6D",X"F9F6FD",X"FAFCF7",X"FFFFFB",X"FEF5F8",X"FEF9FF",X"D4AAE9",X"5D005D",X"C88FD3",X"FFFEFF",X"FFF9FD",X"FAF8FF",X"F8FFFF",X"FBF9FF",X"F0FFF5",X"FFF8FF",X"FFE3FF",X"FF99FF",X"C00695",X"E03DBA",X"AD4594",X"DB87B9",X"C91D97",X"FFDBFF",X"FFFBFF",X"F1F9EE",X"F7F6F1",X"FFF9F7",X"F7FFFF",X"FFC9FA",X"C70096",X"E728B3",X"E6B4E7",X"FFFAFF",X"FFFCFF",X"F6F8F5",X"FFFEF8",X"FCFFFF",X"FFFCF5",X"FFFFFA",X"C3D9D7",X"003130",X"1F5256",X"061E28",X"414449",X"010000",X"756D6B",X"FCFCFA",X"FFFEFF",X"FFFCFF",X"FFFEFF",X"F8FEFC",X"FFFCFF",X"F8DCEA",X"5E4040",X"010100",X"090C15",X"DFD7E6",X"FFFAFC",X"FFFCFF",X"FFFCFF",X"F8FDFF",X"FFFCF5",X"FFFCF9"),
(X"F9FFFF",X"FCFDFF",X"FFF5B8",X"F6DB18",X"F8E203",X"DDD46D",X"F0F3D8",X"FEFFFF",X"FFF9FC",X"FFFCFD",X"FEFCFD",X"FFFDFE",X"FFFDFF",X"FFFDFF",X"FFFCFF",X"FEFEFF",X"FCFEFF",X"91D2FC",X"256DB7",X"000A4F",X"D0BBDA",X"FFFCFD",X"FBFBF9",X"F5F2F9",X"F0FFFF",X"C7FFF8",X"ACE9D7",X"EAFFFF",X"E6FBF4",X"FFFCFD",X"FCF3F8",X"DFFFF9",X"83D7BF",X"00100E",X"000102",X"A6979E",X"FFFAFF",X"FAF9FF",X"FFF2FF",X"FEFCFF",X"FFF2F7",X"FFF8FE",X"FFEFFF",X"FFF8FF",X"E8E4F3",X"828373",X"8C895C",X"BAAD76",X"F7EDE4",X"F4FAF8",X"F5FAF3",X"FFFCFF",X"F7FDF1",X"FFF0FA",X"B058C0",X"75017E",X"410F56",X"CAC8DE",X"FFFBFF",X"F2F2F4",X"EEF9FB",X"EAFFFF",X"C2FFEF",X"B6F0D8",X"EBFFFC",X"FFFDFF",X"F8FFFF",X"F8FFFF",X"C5FFF0",X"15ECA9",X"05CB90",X"45D3AD",X"CFFFFF",X"F8FFFF",X"FAF6F5",X"FDF4F9",X"FFF2FF",X"F1DFFF",X"C489CB",X"E047B1",X"D860B9",X"F9B0E8",X"FFF6FF",X"F8F9F4",X"FFFEF9",X"D5FFFC",X"4EE9BD",X"00CD95",X"A3F1F1",X"F4FFFF",X"FFFEFD",X"F7FFFF",X"F3FDFC",X"F7FFFF",X"FCFAFF",X"FFE1EA",X"D862AC",X"CE056D",X"BE005C",X"FFB8F0",X"FFEFFF",X"F5F5F7",X"F3FFF9",X"EDFFFB",X"FFF8F0",X"817589",X"000500",X"301B00",X"FFE4C1",X"FFFEEF",X"FFF9F0",X"FDF6E4",X"FFFBF4",X"FFFDDF",X"FFF1BA",X"E8E1AB",X"FFFFEF",X"FFF9FF",X"FFFAEA",X"FFF4B9",X"F3C12C",X"DCAD05",X"E8C574",X"FFFBEF",X"F4FFF2",X"FCFDEB",X"FFFFF3",X"FBFEFF",X"E9E8ED",X"EEEDF2",X"FDFDFF",X"F6F6F8",X"FFFFFF",X"FFFFFF",X"FBFBF9",X"FFFFFD",X"FCFFFF",X"F5ECEF",X"FFFFFD",X"F5FEF9",X"FDFBFE",X"FFFFFF",X"DAD1D4",X"57343B",X"811E18",X"A7000E",X"FFB8B9",X"FEFBF6",X"FAFFFF",X"F4FFFA",X"F3FFF1",X"EFFFF8",X"FCFFEC",X"F6FFF1",X"F0FFF4",X"C9ECC4",X"7EAB68",X"608945",X"A1BA93",X"F7FFF8",X"FFFEFF",X"F9FAFC",X"FCFBFF",X"F1FAFF",X"FAEFFF",X"E871B1",X"CE0061",X"D4006A",X"DB65B1",X"FFE6FF",X"FCFEFB",X"F4FFFD",X"FEFEFF",X"E9FEFF",X"A3E4EA",X"D2F3FF",X"FDFDFD",X"FDFDFD",X"FCFCFC",X"FDFDFD",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"F3F7F6",X"FFF7FF",X"FFFBFF",X"F0FFFF",X"95E1FB",X"028FD6",X"0DA4F5",X"299CD2",X"D4F9F2",X"F2FFFF",X"F7FFFD",X"F2FFFF",X"E9FCFF",X"FBFFFF",X"9F99A7",X"D7D4DF",X"FEFDFF",X"FFC1F4",X"B61160",X"9C064D",X"D98DB4",X"FFF3FF",X"FFFDFF",X"FFFBFF",X"E8FDFE",X"FFFEFF",X"FFFBFF",X"FFEFFC",X"A04F7A",X"B0125D",X"960046",X"FF9BD6",X"FFF6FF",X"FFEBF8",X"FDF4F7",X"F3FEFA",X"EAD4E0",X"8C345E",X"820040",X"C94287",X"FFD9F5",X"FFEAFC",X"FFF9FF",X"FFF8FF",X"FFF8FF",X"FFFBFF",X"FFF6FF",X"FEF8FC",X"746A6B",X"010007",X"D6D5E5",X"FFFCFF",X"F3F2F7",X"FBFFFB",X"F1F6F2",X"FFFEFF",X"746578",X"D8CBD2",X"FFF8F1",X"FFFFF3",X"FCFFF4",X"F0F8ED",X"FEFFF4",X"B8B9A7",X"000400",X"000404",X"EDEFEC",X"FFF6ED",X"FFFFFB",X"D2F2FF",X"184B5C",X"001117",X"A1B2AC",X"FFFFFA",X"FFF8FB",X"FFF7FF",X"FFFDFF",X"FFFEFF",X"F1FCF4",X"E2FFF3",X"3DC3C2",X"428F99",X"000717",X"C1BEC7",X"FEFFFF",X"FBFDFA",X"FFFBFF",X"FFF1FB",X"C885D5",X"5C0072",X"C06EC3",X"FFEEF4",X"FFFFF3",X"EDFFF9",X"D9FFF2",X"FFFEFB",X"F1F5F6",X"FFFBFF",X"F2F6F5",X"F7FCFF",X"E1B3D7",X"A22E7F",X"D439B1",X"B30694",X"BE2E9F",X"FED9FF",X"FFFDFF",X"FEFFFA",X"FFFFF8",X"FEFBF4",X"FCFFFF",X"FFC8FB",X"DA00B5",X"BF058E",X"DF92BE",X"FAF9F4",X"FFF3FC",X"F7FFF8",X"F4FFED",X"F1FFF6",X"FAFFF4",X"FCFFFB",X"FAF5FC",X"DBD3E8",X"0C1222",X"000307",X"301F18",X"280000",X"9F7078",X"FFFAFB",X"FAFEFD",X"F6F4F5",X"FFF5F6",X"FFFFFD",X"FCFFFF",X"CDCED3",X"251F29",X"000D24",X"000325",X"D2D4E9",X"FEFFFA",X"ECFDEB",X"F4FFF7",X"FFFFFA",X"EFF0E0",X"F5EEE4"),
(X"F7FEFF",X"FAFBFF",X"FCEEB1",X"E8CD0A",X"F1DB00",X"EEE57E",X"FDFFE5",X"FAFBFF",X"FFF9FC",X"FFFBFC",X"FEFCFD",X"FFFDFE",X"FFFDFF",X"FFFDFF",X"FFFDFF",X"FEFEFF",X"F5F7FF",X"80C1EB",X"2D75BF",X"071156",X"A994B3",X"FFF8F9",X"FFFFFD",X"FCF9FF",X"E0F6F4",X"BEFFEF",X"4A8775",X"D5F5EA",X"F1FFFF",X"FDF9FA",X"FFF6FB",X"DEFFF8",X"7FD3BB",X"000604",X"000102",X"97888F",X"FEF1FA",X"FEFDFF",X"FFF4FF",X"F8F6FF",X"FFFAFF",X"FFF8FE",X"FFF7FF",X"DDCFE9",X"595564",X"0B0C00",X"070400",X"E5D8A1",X"FFFCF3",X"FBFFFF",X"F8FDF6",X"F9F6FF",X"F9FFF3",X"FFF3FD",X"AF57BF",X"76027F",X"320047",X"C8C6DC",X"FFFBFF",X"FFFFFF",X"F0FBFD",X"DBFBF0",X"95E2C2",X"70AA92",X"E6FDF7",X"FFFDFF",X"F3FEFA",X"F4FEFD",X"C0FDEB",X"00D18E",X"13D99E",X"46D4AE",X"BEF5F0",X"EEF8FA",X"FFFDFC",X"FFFCFF",X"FFEDFF",X"FFF5FF",X"FFCDFF",X"F55CC6",X"D961BA",X"843B73",X"B4A6B5",X"FBFCF7",X"FFFFFA",X"B6F1DD",X"16B185",X"1AE7AF",X"B2FFFF",X"F1FFFE",X"FDF9F8",X"F8FFFF",X"F8FFFF",X"F8FFFF",X"FBF9FF",X"FFF4FD",X"FD87D1",X"CA0169",X"CE0A6C",X"CE6FA7",X"F4DDF1",X"FFFFFF",X"F0FFF6",X"EDFFFB",X"F3ECE4",X"4F4357",X"000800",X"978253",X"FFE1BE",X"FFFFF0",X"FDF4EB",X"FFFEEC",X"FFF6EF",X"FFF5D7",X"D0C18A",X"DED7A1",X"FFFFEF",X"F9F1FC",X"FFFCEC",X"EDDEA3",X"E9B722",X"E1B20A",X"EDCA79",X"FFFFF3",X"F4FFF2",X"F7F8E6",X"FFFFF3",X"F2F5FF",X"6E6D72",X"C8C7CC",X"FCFCFE",X"FBFBFD",X"FFFFFF",X"FCFCFC",X"FFFFFD",X"FEFEFC",X"F8FCFF",X"FFFCFF",X"FEFEFC",X"F0F9F4",X"F8F6F9",X"FFFFFF",X"DBD2D5",X"1E0002",X"801D17",X"A8000F",X"FFADAE",X"FCF9F4",X"F5FBFB",X"F4FFFA",X"EBF7E9",X"EDFFF6",X"F6FEE6",X"EAF5E5",X"B8CDBC",X"71946C",X"5C8946",X"99C27E",X"DFF8D1",X"F6FFF7",X"FCFAFF",X"FEFFFF",X"FFFEFF",X"F8FFFF",X"FBF0FF",X"D05999",X"D60269",X"D4006A",X"D45EAA",X"FFDDFE",X"FEFFFD",X"E4F5ED",X"FEFEFF",X"D6EBFE",X"226369",X"AECFDE",X"FCFCFC",X"FCFCFC",X"FCFCFC",X"FDFDFD",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FCFFFF",X"FFF8FF",X"FDF7FF",X"E8FDFF",X"7FCBE5",X"0794DB",X"0FA6F7",X"2C9FD5",X"D7FCF5",X"F0FFFD",X"F6FFFC",X"E8FBF9",X"E4F7FB",X"D6DAE6",X"06000E",X"D2CFDA",X"FCFBFF",X"DE84B7",X"AA0554",X"AB155C",X"FFC5EC",X"FFF7FF",X"FFFBFF",X"FFFDFF",X"F0FFFF",X"FEFDFF",X"FFFBFF",X"FDEDFA",X"E392BD",X"A2044F",X"B31663",X"B14984",X"F2DAE8",X"FFF6FF",X"FFF7FA",X"F8FFFF",X"FFF6FF",X"D880AA",X"910F4F",X"940D52",X"C28DA9",X"FFE7F9",X"FFF2FC",X"FFFAFF",X"FFFBFF",X"FDF3FE",X"F6ECF5",X"AEA8AC",X"0A0001",X"84818A",X"F9F8FF",X"FDF9FF",X"FEFDFF",X"F9FFF9",X"F8FDF9",X"FCFAFF",X"897A8D",X"4F4249",X"FCF3EC",X"F6F7E9",X"F9FFF1",X"F6FEF3",X"F9FDEF",X"80816F",X"000400",X"A5B1B1",X"F9FBF8",X"FFF4EB",X"FDFCF8",X"A2C2CF",X"285B6C",X"57868C",X"E6F7F1",X"FFFFFA",X"FFF5F8",X"FFFAFF",X"FDFBFF",X"FFFEFF",X"F6FFF9",X"E6FFF7",X"75FBFA",X"226F79",X"021323",X"5E5B64",X"F2F4F3",X"FBFDFA",X"FFF9FE",X"FEEDF7",X"AF6CBC",X"6A0680",X"903E93",X"FFE9EF",X"FEFAEE",X"EEFFFA",X"E4FFFD",X"FDF8F5",X"FCFFFF",X"FFFDFF",X"F9FDFC",X"FAFFFF",X"FFDFFF",X"FF93E4",X"CE33AB",X"E93CCA",X"CA3AAB",X"FFDCFF",X"FCFAFD",X"FBFEF7",X"FBF8F1",X"F9F6EF",X"FCFFFF",X"FFC5F8",X"D600B1",X"F43AC3",X"BF729E",X"FBFAF5",X"FFF8FF",X"EDFBEE",X"F4FFED",X"F5FFFA",X"FCFFF6",X"F6FBF5",X"FFFDFF",X"FFF9FF",X"BDC3D3",X"000509",X"200F08",X"450F05",X"AB7C84",X"FFF5F6",X"F9FDFC",X"FFFEFF",X"FFFAFB",X"F1F0EE",X"F7FBFC",X"C3C4C9",X"030007",X"32485F",X"2E4668",X"C3C5DA",X"FEFFFA",X"F1FFF0",X"F4FFF7",X"FBFAF5",X"A4A595",X"D7D0C6"),
(X"FBFFF4",X"F8FAED",X"F8F898",X"EBE52B",X"DDD228",X"E6E863",X"FAFEC3",X"FFFFF3",X"FFF8F9",X"FFFBFA",X"FDFDFD",X"FFFDFF",X"FFFCFF",X"FFFCFF",X"FEFEFF",X"FBFFFF",X"FAEAF5",X"567091",X"356B97",X"153355",X"00101D",X"66A094",X"9CFFE4",X"9FFFE6",X"86FCDA",X"4ACEA6",X"7BCBB2",X"E8F7F2",X"FAFAFA",X"FFF1F8",X"FFF8FF",X"D9FFFA",X"70DCBC",X"21604F",X"000704",X"070002",X"AB97A3",X"FED8F1",X"FFC4E8",X"FFCCF3",X"FFBCFF",X"F3ACF2",X"A961AA",X"4A105C",X"1A002F",X"716279",X"E3D9E1",X"FFFBFF",X"F5FFFE",X"E7F9E9",X"FBFFFA",X"F7F9F8",X"FFFFFA",X"E6C1E0",X"621269",X"661572",X"33002D",X"435257",X"6D7170",X"70CAB1",X"7EFFDB",X"75E5BD",X"14AB76",X"94E7D5",X"F2FFFE",X"FFF8FE",X"FCF8F9",X"FDFFFE",X"C6F6E6",X"20CC94",X"29D09C",X"0FC28B",X"88F0D5",X"E7FFFF",X"FBFFFD",X"E9F9EF",X"FFFCFD",X"FFFBFA",X"F1F3E8",X"EAD6CF",X"B47EB2",X"784E72",X"010005",X"84A296",X"C3FFEA",X"5FDCB4",X"17C48F",X"36E0AF",X"D1EFF9",X"FFFDFF",X"FFF8FF",X"FFFCFF",X"FFFDF1",X"FFFAF8",X"FBF8FF",X"FCFBF9",X"EFC3E6",X"A61560",X"CC0A6A",X"9A024F",X"FFA7D6",X"FFE6FA",X"FFF2F8",X"FFF5FA",X"F5E9EB",X"080122",X"1D1500",X"CEAD42",X"E9CD5F",X"FBF7AE",X"EFE6A1",X"FFF093",X"ECE16D",X"E1CE67",X"B89F4D",X"EED9AC",X"FFFBFA",X"FFF7FF",X"FFFBEA",X"F1DA96",X"D7BA21",X"D6C106",X"D3BC38",X"F7E498",X"FFF2A7",X"FFF38F",X"E6D06D",X"91704D",X"060606",X"C7C7C7",X"FFFFFF",X"FAFAFC",X"FFFFFF",X"FEFEFF",X"FCFCFC",X"FFFFFF",X"F9FFFF",X"FFF8FC",X"FBF7F6",X"FBFFFD",X"FFFEFF",X"FEFFFF",X"ADB2B5",X"070002",X"362720",X"862933",X"B25C69",X"977D88",X"7B8386",X"A5C1AB",X"C4E6C5",X"A8C6AA",X"9AB081",X"8CA17A",X"718667",X"6C8462",X"9DB790",X"E3F6DA",X"FCFFFB",X"FEF6FF",X"FBFFFF",X"FAFAFA",X"F3F3F1",X"FCFFFF",X"FFE6FA",X"AF447A",X"B00D5C",X"AC0356",X"B01D75",X"CB6DA2",X"9D7389",X"9FB0B8",X"82ABBD",X"68A4BE",X"519AAB",X"CFE7FF",X"FCFCFC",X"FCFCFC",X"FCFCFC",X"FDFDFD",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"F7FBED",X"EEF9FD",X"F8FFFF",X"E0FCFF",X"6BB8D4",X"2495CD",X"168ECA",X"108EBE",X"6ED5FE",X"A7F8FF",X"AAEBFF",X"AEF0FF",X"90C6E2",X"3F546F",X"000010",X"E4DAE5",X"FFB9E0",X"96064B",X"BF0559",X"A51A5D",X"FAC5E3",X"FFFEFF",X"FFFFFF",X"FFF3FB",X"FFF6FF",X"FFF8FE",X"F3FFFF",X"F2FFFF",X"FDCCEC",X"A01358",X"B10557",X"A00E55",X"E489B5",X"FFEAFA",X"F7FDFB",X"F7F1F1",X"FFF8FF",X"F6E4F2",X"A9698B",X"880B43",X"980442",X"F67EAE",X"FFC0E6",X"FFC2E7",X"FFB5E2",X"FFBCE7",X"CB88A7",X"190005",X"6B666C",X"FBF2F7",X"FEF9FD",X"FAFEFD",X"FBFFFF",X"FCFAFD",X"FDF8FC",X"FFFFFF",X"71867F",X"000C00",X"979656",X"FFFF9E",X"FFFF8A",X"FFFA8A",X"D6C870",X"8E813D",X"A79686",X"F7EDE3",X"FBFFFE",X"ECFFFF",X"B9F2FF",X"4AA6BD",X"30A3B8",X"33AEBE",X"C4FCFD",X"EDFFFF",X"FFFDFC",X"FFFFF1",X"FBFEEB",X"FFFEF8",X"FFFAF9",X"FFF9F1",X"C7FFFF",X"609094",X"041C20",X"000004",X"99979A",X"FEFFFF",X"FEF7FF",X"FFF0FF",X"8D3486",X"460C70",X"630367",X"E3C0EA",X"F4FFFF",X"FFF6FF",X"F5F4EF",X"FFF2F6",X"FFFFF4",X"EBEFEE",X"FCF4FF",X"FFF9FF",X"F6FCFA",X"FFFEFF",X"E2A6D9",X"C852B0",X"A85293",X"F0DDF3",X"F4FDFC",X"FCFCFE",X"FFF9FC",X"FFFFFB",X"FCF7FD",X"E4B2D8",X"99146F",X"92557F",X"471016",X"E2D0CC",X"F8FEFF",X"FCFFFF",X"FFF7FA",X"F7F4FF",X"F8FFFF",X"FCFFFF",X"FDF4F9",X"FDF3FC",X"F3F2F7",X"C7BBBD",X"500911",X"880316",X"AC797E",X"FFF4F5",X"F0F9F8",X"FCFDFF",X"FEF9F6",X"FCFDF8",X"F9FFFF",X"ACB3BB",X"000A14",X"398A9D",X"3D9AA9",X"4C7179",X"898083",X"969792",X"A5A89F",X"A58C88",X"6B6350",X"E2D6C8"),
(X"F7FFF0",X"CFD1C4",X"CBCB6B",X"EDE72D",X"E4D92F",X"DBDD58",X"CCD095",X"CDCEC0",X"FFF9FA",X"FFFBFA",X"FDFDFD",X"FFFDFF",X"FFFCFF",X"FFFCFF",X"FEFEFF",X"FBFFFF",X"9E8E99",X"001536",X"3E74A0",X"375577",X"20303D",X"1B5549",X"5BBFA3",X"4EB395",X"43B997",X"199D75",X"95E5CC",X"F5FFFF",X"FCFCFC",X"FFF1F8",X"FFFAFF",X"94C2B5",X"54C0A0",X"6DAC9B",X"000603",X"11060C",X"0D0005",X"27011A",X"4A0E32",X"470F36",X"44004B",X"520B51",X"570F58",X"9B61AD",X"CDAAE2",X"F4E5FC",X"FFFBFF",X"FFFAFF",X"F6FFFF",X"F1FFF3",X"EEF5ED",X"FEFFFF",X"F6F7F1",X"9F7A99",X"722279",X"863592",X"6C3866",X"253439",X"080C0B",X"217B62",X"3FC39C",X"40B088",X"17AE79",X"AAFDEB",X"EFFEFB",X"FFF9FF",X"FFFEFF",X"F0F2F1",X"96C6B6",X"22CE96",X"30D7A3",X"39ECB5",X"61C9AE",X"9BB8B3",X"E8EEEA",X"F0FFF6",X"FFF8F9",X"FFFBFA",X"FDFFF4",X"FFF2EB",X"FAC4F8",X"956B8F",X"39363D",X"224034",X"6AA891",X"3AB78F",X"38E5B0",X"22CC9B",X"ABC9D3",X"F9F4FA",X"FFF8FF",X"FFF9FF",X"FFFBEF",X"FFFDFB",X"FFFDFF",X"F7F6F4",X"FFE0FF",X"D4438E",X"D91777",X"CC3481",X"953867",X"C297AB",X"F7E6EC",X"FFF3F8",X"A29698",X"2B2445",X"776F5A",X"D8B74C",X"D6BA4C",X"B2AE65",X"B3AA65",X"B7A84B",X"B2A733",X"AA9730",X"BCA351",X"FEE9BC",X"FFF9F8",X"FFF2FF",X"E5D2C1",X"CFB874",X"DDC027",X"E1CC11",X"C9B22E",X"C5B266",X"B5A55A",X"BAA844",X"BBA542",X"8C6B48",X"696969",X"EBEBEB",X"FDFDFF",X"FAFAFC",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FDFDFD",X"F6FEFF",X"FFFBFF",X"FFFEFD",X"F1F7F3",X"FFFEFF",X"D5D6DB",X"33383B",X"21161C",X"0C0000",X"5C0009",X"4E0005",X"110002",X"000205",X"4F6B55",X"789A79",X"567458",X"778D5E",X"80956E",X"98AD8E",X"C6DEBC",X"EEFFE1",X"F5FFEC",X"F5FAF4",X"FFF8FF",X"F3F8FB",X"FFFFFF",X"FFFFFD",X"FAFEFF",X"DDC0D4",X"A1366C",X"C92675",X"D93083",X"C43189",X"83255A",X"1C0008",X"00050D",X"133C4E",X"3E7A94",X"6FB8C9",X"E7FFFF",X"FDFDFD",X"FDFDFD",X"FCFCFC",X"FDFDFD",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFFF4",X"F7FFFF",X"F8FFFF",X"C1DDE0",X"519EBA",X"2D9ED6",X"29A1DD",X"2CAADA",X"2D94BD",X"3586B1",X"3879A1",X"327494",X"5A90AC",X"1A2F4A",X"9B98AB",X"D0C6D1",X"883D64",X"B8286D",X"E92F83",X"AA1F62",X"AF7A98",X"EBEAEF",X"FAFAFC",X"FFF9FF",X"FFF2FD",X"FFFBFF",X"F5FFFF",X"EEFFFF",X"FFDDFD",X"E4579C",X"B70B5D",X"C5337A",X"872C58",X"B192A2",X"E2E8E6",X"FFF9F9",X"FFF6FE",X"FFF8FF",X"FFCFF1",X"FF92CA",X"BB2765",X"7E0636",X"6C0C32",X"701439",X"821B48",X"6B0A35",X"5A1736",X"B08B9C",X"FFFDFF",X"FEF5FA",X"FBF6FA",X"FCFFFF",X"F0F6F6",X"FFFEFF",X"F8F3F7",X"FFFFFF",X"8A9F98",X"000900",X"696828",X"B0A644",X"B7A833",X"B3A636",X"B9AB53",X"D7CA86",X"FFF2E2",X"FFFDF3",X"EFF3F2",X"C8E1E8",X"619AAB",X"429EB5",X"3EB1C6",X"2FAABA",X"96CECF",X"E3F6FD",X"FFFEFD",X"FFFFF0",X"FEFFEE",X"FFFDF7",X"FFF7F6",X"FFFEF6",X"C3FEFF",X"82B2B6",X"3E565A",X"3F4044",X"050306",X"8F9092",X"E8E1E9",X"BFAAB9",X"7A2173",X"8349AD",X"88288C",X"83608A",X"B6C4CF",X"FFF2FD",X"FFFFFA",X"FFF7FB",X"FDF9EE",X"FCFFFF",X"FFFBFF",X"FCEEFB",X"F7FDFB",X"F4F3F9",X"FFE3FF",X"FFA5FF",X"9F498A",X"F2DFF5",X"F9FFFF",X"F7F7F9",X"F9F0F3",X"FFFFFB",X"D0CBD1",X"825076",X"BC3792",X"672A54",X"4B141A",X"65534F",X"E9EFFD",X"F6F9FF",X"FFF2F5",X"FFFCFF",X"F8FFFF",X"F5F9FA",X"FFFCFF",X"FFFBFF",X"FCFBFF",X"FFF3F5",X"F6AFB7",X"890417",X"C39095",X"FFF7F8",X"F3FCFB",X"F8F9FB",X"FFFBF8",X"FEFFFA",X"E5EEED",X"737A82",X"466872",X"62B3C6",X"46A3B2",X"668B93",X"0B0205",X"070803",X"000200",X"523935",X"7E7663",X"E9DDCF"),
(X"FFF3FF",X"F7EFED",X"F5F5DD",X"FBFEDF",X"F4F2E5",X"FFFFCA",X"FAEBE4",X"FBE6EB",X"FFFCFB",X"FDFDFB",X"FDFFFE",X"FDFEFF",X"FFFEFF",X"FEFEFF",X"FBFFFF",X"F8FFFF",X"E7F4E3",X"EAEEF1",X"EFF8FD",X"F6F2F1",X"FFEBEF",X"EFF4F7",X"C7E8E1",X"E0F2E6",X"D9EBEB",X"C8FAEE",X"EEFFFF",X"FDFBFC",X"F1FFFB",X"FFFEFF",X"FFF6FD",X"DAF8F0",X"E5F5F4",X"D5F4EC",X"C9C4C8",X"A8A7AC",X"AAAAB2",X"C1A1B9",X"BDA0BE",X"B499BA",X"B4ABBE",X"D2C0CE",X"FFE9F6",X"FFE6F9",X"FFFAFF",X"FFFEFF",X"FEFEFC",X"FCFAFB",X"FFFAF0",X"FFF9FF",X"FFF7FF",X"FFFFF4",X"F2F5FC",X"F7DAFF",X"FFE0F5",X"FBEFF9",X"FAEEFA",X"F0EFED",X"F5DEE4",X"DAE8EB",X"CEEEE9",X"E8FCF3",X"D2F3EC",X"F6F7FF",X"F5FFFF",X"FFF6FD",X"F8F8F8",X"FBFDFA",X"DDF2E9",X"E4F9F2",X"CAFAEC",X"D4F9F1",X"DEF7FE",X"D7E7E7",X"FFFFFB",X"FFFFF8",X"F6FDF6",X"F2FFFF",X"F5F9FF",X"FFF8FF",X"FFF1FF",X"F9E9F6",X"FAEDF6",X"F2FBFA",X"D9FEF7",X"E6FFFF",X"E1EBED",X"DCF7F0",X"D8F5E3",X"F4FCE7",X"FFFCFE",X"FCFFFF",X"F9FFFB",X"F6F7FC",X"FEFEFF",X"F9FFF1",X"F8F7FC",X"FCE9FD",X"F6E8FF",X"E7DDF8",X"F8E6FE",X"E7E4EF",X"F8FFFF",X"F3F1F2",X"E3F3E8",X"E9F2F7",X"FFE7E0",X"FFFEDD",X"EDFBE2",X"F1F2E0",X"F5F0D3",X"F4E7D6",X"F5F1D6",X"E7DAD1",X"F3E3E3",X"FFFFF4",X"F6FFF7",X"F4FFFF",X"EFF6EF",X"F3EEDB",X"F7F3E7",X"F8FAD2",X"F9F6D5",X"FFF9DE",X"F4EBDC",X"EFECDB",X"ECF0CF",X"E9E8E4",X"F7F7F5",X"FFFFFF",X"F9F9F9",X"FDFDFF",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"F9F9FB",X"F8FFFF",X"FFF9FD",X"FFFAF7",X"F7FDFB",X"FAF8FD",X"F5F8FF",X"E2F0F3",X"DEE2E5",X"BEB1C2",X"AFA3A3",X"ABA6A3",X"9D9DA9",X"A09AA4",X"C3C6B5",X"B2CBA4",X"B8CCA9",X"C5E3CB",X"E1F7E2",X"F7FFF5",X"F9FFF9",X"F8FCFD",X"FEFDFF",X"FFFCFF",X"FFFBFF",X"FFFFFF",X"FFFBFD",X"FFFAF7",X"FAFCF7",X"FDF2FA",X"F3D6EC",X"F7DDF6",X"ECDFF3",X"FCE2EF",X"ECEDE7",X"F1E2DB",X"E7E7E9",X"DBEEFD",X"DEE2FF",X"EAF1FF",X"F4FFFF",X"FEFEFE",X"FDFDFD",X"FDFDFD",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFF8F4",X"F5FCFF",X"FFFCFD",X"FAE8E4",X"D9E5F1",X"DEF4FF",X"E6F9FD",X"D2FAFA",X"DFF9F6",X"EDF8FA",X"DFECF2",X"D0EDF1",X"CCEDF2",X"E2F1F8",X"F3F1F4",X"F0EBE7",X"F2E4F3",X"EFEBFA",X"E9E0F5",X"F5DBF4",X"F9E1F1",X"FBF7F8",X"F8FFFB",X"F6FFF8",X"FEFFFD",X"F2F9F2",X"FEFFFB",X"FFF9FE",X"FFF4FF",X"F7F2FF",X"EBDDF6",X"FFE4FF",X"F7E9FF",X"ECDAEA",X"FAEFF3",X"F9FFFA",X"F7FFFA",X"FAF6F7",X"FFFBFF",X"FBF5F9",X"FFEBFF",X"D1BACC",X"BC9DAF",X"C298AE",X"BE90AC",X"D0ADC5",X"F4E3F3",X"F7F8FD",X"F1F4FB",X"FFFCFD",X"FFFDF4",X"F7FFF7",X"F7FFFE",X"FFFBFF",X"FFFBFF",X"FBFDFA",X"FEE7F9",X"ABA7A4",X"A9B59D",X"CED5B4",X"D0C2A8",X"D8BFAB",X"F5E7CD",X"FFFFE0",X"FFFCFF",X"FFF6F7",X"FFFEFB",X"DAEFF2",X"CDF0F2",X"E1FFFA",X"DFFEF6",X"CEF8F6",X"DEE9E5",X"FFF9FF",X"FFF9FF",X"F2FCF3",X"F7FFFF",X"FCFDFF",X"FFFBFF",X"FFFCFF",X"FFF8FF",X"EFF9FA",X"E3F8F3",X"F2F8F6",X"F5EFF3",X"FAF7FE",X"F0EDF8",X"F4E3F5",X"FBE4EC",X"EAE5FC",X"F6E4FE",X"F6E3F6",X"F5E9F7",X"FFF6F7",X"FFFFFA",X"EFFBFF",X"FFFDFF",X"EDF7F9",X"FFFDFF",X"FFF9FD",X"FFFFFF",X"FFFBFF",X"FFFBFB",X"EAFFF3",X"FFD9F0",X"FFF9F9",X"ECFDF5",X"FFFDFF",X"FFFAFF",X"FBFFFE",X"FBEEF5",X"FFDBF6",X"FCDFF1",X"E3F4EE",X"FFF3F0",X"EAE7F2",X"EEF2FF",X"FFFAFF",X"FEFFEF",X"FDFAF5",X"FFFAFF",X"FFFBFF",X"FAF9F4",X"EEFCEF",X"F5FFF6",X"FFFBFB",X"FFEEF1",X"F6E6E6",X"FAE6DF",X"FFFFFA",X"F9FDFE",X"FEFFFF",X"FEFFFB",X"F2FEF4",X"FCFDFF",X"F2E0F0",X"E7F4ED",X"EAF1FF",X"E6F6FF",X"EDFEF6",X"E2E7E3",X"E5EDF0",X"E5EBE9",X"EEDBD5",X"EEE0D3",X"FFFCF4"),
(X"FFF9FF",X"FFFDFB",X"FEFEE6",X"FDFFE1",X"FFFEF1",X"FFFFCD",X"FFF4ED",X"FFF8FD",X"FFFDFC",X"FEFEFC",X"FEFFFF",X"FEFFFF",X"FFFEFF",X"FFFFFF",X"FBFFFF",X"F8FFFF",X"F7FFF3",X"FCFFFF",X"F8FFFF",X"FFFCFB",X"FFF7FB",X"F6FBFE",X"E9FFFF",X"F4FFFA",X"F2FFFF",X"D9FFFF",X"ECFFFF",X"FFFEFF",X"F4FFFE",X"FFFDFE",X"FFFAFF",X"EAFFFF",X"F1FFFF",X"EAFFFF",X"FEF9FD",X"FFFEFF",X"F9F9FF",X"FFEFFF",X"FFF3FF",X"FFF3FF",X"FFFAFF",X"FFF8FF",X"FFEEFB",X"FFF5FF",X"FFF5FF",X"FDFBFE",X"FDFDFB",X"FFFEFF",X"FFFEF4",X"FFFAFF",X"FFF6FF",X"FFFFF4",X"FCFFFF",X"FFF1FF",X"FFF1FF",X"FFFAFF",X"FFF7FF",X"FFFFFD",X"FFF3F9",X"F5FFFF",X"E9FFFF",X"E9FDF4",X"E9FFFF",X"FCFDFF",X"F1FFFF",X"FFFAFF",X"FCFCFC",X"FDFFFC",X"F0FFFC",X"EBFFF9",X"DFFFFF",X"E6FFFF",X"ECFFFF",X"F4FFFF",X"F9FAF5",X"FFFFF8",X"F8FFF8",X"F4FFFF",X"FBFFFF",X"FFF7FF",X"FFF7FF",X"FFF9FF",X"FFF5FE",X"F9FFFF",X"E6FFFF",X"E7FFFF",X"F8FFFF",X"EDFFFF",X"EDFFF8",X"F8FFEB",X"FFFDFF",X"FAFDFF",X"F9FFFB",X"FEFFFF",X"FEFEFF",X"F7FFEF",X"FFFEFF",X"FFF3FF",X"FFF8FF",X"FFF9FF",X"FFF4FF",X"FEFBFF",X"F8FFFF",X"FFFEFF",X"F4FFF9",X"F8FFFF",X"FFF8F1",X"FFFFDF",X"F7FFEC",X"FFFFEF",X"FFFFE4",X"FFF9E8",X"FFFFE6",X"FFFBF2",X"FFFAFA",X"FFFFF4",X"F4FFF5",X"F2FFFF",X"FBFFFB",X"FFFFEC",X"FFFFF3",X"FFFFDA",X"FFFFE1",X"FFFFE4",X"FFF7E8",X"FFFFEF",X"FAFEDD",X"FFFFFB",X"FEFEFC",X"FCFCFC",X"FFFFFF",X"FDFDFF",X"FFFFFF",X"FCFCFE",X"FFFFFF",X"FFFFFF",X"F6FFFF",X"FFFBFF",X"FFFEFB",X"FBFFFF",X"FFFEFF",X"F8FBFF",X"F5FFFF",X"F8FCFF",X"FFF9FF",X"FFF9F9",X"FFFAF7",X"FEFEFF",X"FFFCFF",X"FFFFF1",X"F0FFE2",X"F5FFE6",X"EDFFF3",X"EEFFEF",X"F6FFF4",X"FBFFFB",X"FCFFFF",X"FEFDFF",X"FFFCFF",X"FFF9FF",X"FFFFFF",X"FFF4F6",X"FFFDFA",X"FEFFFB",X"FFFAFF",X"FFF4FF",X"FFF2FF",X"FFF9FF",X"FFF6FF",X"FFFFFA",X"FFFAF3",X"FEFEFF",X"EEFFFF",X"F9FDFF",X"F5FCFF",X"F6FFFF",X"FFFFFF",X"FEFEFE",X"FEFEFE",X"FEFEFE",X"FFFFFF",X"FFFFFF",X"FFFFFF",X"FEFEFE",X"FFFAF6",X"F7FEFF",X"FFFCFD",X"FFF8F4",X"F5FFFF",X"EAFFFF",X"F1FFFF",X"DEFFFF",X"EDFFFF",X"F4FFFF",X"F5FFFF",X"EAFFFF",X"E7FFFF",X"F4FFFF",X"FFFEFF",X"FFFEFA",X"FFF6FF",X"FFFCFF",X"FFFAFF",X"FFF3FF",X"FFF3FF",X"FFFEFF",X"F8FFFB",X"F8FFFA",X"FEFFFD",X"FBFFFB",X"F9FBF6",X"FFFCFF",X"FFF7FF",X"FEF9FF",X"FFF8FF",X"FFF0FF",X"FFF8FF",X"FFF5FF",X"FFFBFF",X"F9FFFA",X"F7FFFA",X"FFFEFF",X"FFFBFF",X"FFFBFF",X"FFF0FF",X"FFF6FF",X"FFEFFF",X"FFEFFF",X"FFEEFF",X"FFECFF",X"FFF6FF",X"FEFFFF",X"FCFFFF",X"FFFBFC",X"FEFAF1",X"F8FFF8",X"F7FFFE",X"FFF9FF",X"FFFAFF",X"FDFFFC",X"FFF6FF",X"FFFBF8",X"F5FFE9",X"FEFFE4",X"FFFEE4",X"FFFAE6",X"FFFDE3",X"FFFFE1",X"FCF9FF",X"FFFCFD",X"FFFCF9",X"F0FFFF",X"E6FFFF",X"E3FFFC",X"EAFFFF",X"E2FFFF",X"F8FFFF",X"FFF5FF",X"FFF8FF",X"F9FFFA",X"F7FFFF",X"F4F5FF",X"FFFBFF",X"FFFCFF",X"FFF5FF",X"F8FFFF",X"F1FFFF",X"FBFFFF",X"FAF4F8",X"FCF9FF",X"FFFCFF",X"FFF8FF",X"FFF7FF",X"FFFBFF",X"FFF3FF",X"FFF7FF",X"FFF6FF",X"FFFAFB",X"FFFFFA",X"F5FFFF",X"FFFDFF",X"F8FFFF",X"FDF8FC",X"FFFBFF",X"FFFFFF",X"FFF7FB",X"FFFAFA",X"F0FFF9",X"FFEEFF",X"FFFDFD",X"F3FFFC",X"FFFDFF",X"FFF9FF",X"FCFFFF",X"FFF5FC",X"FFF0FF",X"FFF4FF",X"F4FFFF",X"FFF5F2",X"FFFDFF",X"F9FDFF",X"FFFAFF",X"F2F7E3",X"FFFFFA",X"FFFDFF",X"FFFBFF",X"FFFFFA",X"F7FFF8",X"F9FFFA",X"FFFAFA",X"FFF8FB",X"FFF7F7",X"FFFAF3",X"FFFCF7",X"FCFFFF",X"FBFCFE",X"FBFDF8",X"F8FFFA",X"FCFDFF",X"FFF8FF",X"F7FFFD",X"F8FFFF",X"EBFBFF",X"F4FFFD",X"FCFFFD",X"F4FCFF",X"FBFFFF",X"FFF8F2",X"FFFCEF",X"FFF9F1")
);
begin
   -- addr register to infer block RAM
   process (clock)
   begin
      if (rising_edge(clock)) then
        if ((unsigned(frst_pixel_v)-1 < unsigned(line_data)) and (unsigned(line_data) < X"A0"+unsigned(frst_pixel_v))
            and (unsigned(frst_pixel_h)-1 < unsigned(column_data)) and (unsigned(column_data) < X"14A"+unsigned(frst_pixel_h))) then -- 330 / 160
          tx <= ROM(to_integer(unsigned(line_data)-unsigned(frst_pixel_v)), to_integer(unsigned(column_data)-unsigned(frst_pixel_h)));
        
        else
          tx <= (others=>'1');
        end if;
      end if;
   end process;

   data <= tx;
end Behavioral;